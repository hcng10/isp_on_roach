//
module ComputeBgNoise(
    input fifodata,
    input periodcount,
    output 
);
endmodule
