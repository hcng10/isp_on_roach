//this module implement the data memory
//use this memory to store the detected object
//for further processing 
