module ROM (addr,data);
input [12:0] addr;
output reg signed [31:0] data;
always@(*)
case(addr)
1: data <= 32'Hffffffed;
2: data <= 32'Hffffffef;
3: data <= 32'Hffffffea;
4: data <= 32'Hffffffe9;
5: data <= 32'Hffffffeb;
6: data <= 32'Hffffffeb;
7: data <= 32'Hfffffff0;
8: data <= 32'Hffffffe6;
9: data <= 32'Hffffffea;
10: data <= 32'Hfffffff0;
11: data <= 32'Hffffffec;
12: data <= 32'Hfffffff0;
13: data <= 32'Hfffffff1;
14: data <= 32'Hffffffef;
15: data <= 32'Hfffffff4;
16: data <= 32'Hfffffff4;
17: data <= 32'Hfffffff2;
18: data <= 32'Hfffffff4;
19: data <= 32'Hfffffff7;
20: data <= 32'Hfffffff2;
21: data <= 32'Hfffffff7;
22: data <= 32'Hfffffff5;
23: data <= 32'Hfffffff4;
24: data <= 32'Hfffffff2;
25: data <= 32'Hfffffffa;
26: data <= 32'Hfffffff4;
27: data <= 32'Hfffffff5;
28: data <= 32'Hfffffff8;
29: data <= 32'Hfffffff5;
30: data <= 32'Hfffffff5;
31: data <= 32'Hfffffff4;
32: data <= 32'Hfffffff4;
33: data <= 32'Hfffffff8;
34: data <= 32'Hfffffff3;
35: data <= 32'Hfffffff1;
36: data <= 32'Hfffffff6;
37: data <= 32'Hfffffff2;
38: data <= 32'Hfffffff3;
39: data <= 32'Hfffffff4;
40: data <= 32'Hfffffff0;
41: data <= 32'Hfffffff0;
42: data <= 32'Hfffffff4;
43: data <= 32'Hfffffff2;
44: data <= 32'Hfffffff3;
45: data <= 32'Hfffffff4;
46: data <= 32'Hfffffff2;
47: data <= 32'Hfffffff4;
48: data <= 32'Hfffffff5;
49: data <= 32'Hfffffff0;
50: data <= 32'Hfffffff8;
51: data <= 32'Hfffffff2;
52: data <= 32'Hfffffff8;
53: data <= 32'Hfffffff7;
54: data <= 32'Hfffffff5;
55: data <= 32'Hfffffff5;
56: data <= 32'Hfffffff9;
57: data <= 32'Hfffffff5;
58: data <= 32'Hfffffff3;
59: data <= 32'Hfffffff6;
60: data <= 32'Hfffffff5;
61: data <= 32'Hfffffff6;
62: data <= 32'Hfffffff2;
63: data <= 32'Hfffffff5;
64: data <= 32'Hfffffff3;
65: data <= 32'Hffffffef;
66: data <= 32'Hfffffff4;
67: data <= 32'Hfffffff5;
68: data <= 32'Hfffffff0;
69: data <= 32'Hfffffff6;
70: data <= 32'Hfffffff7;
71: data <= 32'Hfffffff2;
72: data <= 32'Hfffffff7;
73: data <= 32'Hfffffff4;
74: data <= 32'Hfffffff6;
75: data <= 32'Hfffffff1;
76: data <= 32'Hfffffff3;
77: data <= 32'Hfffffff7;
78: data <= 32'Hfffffff2;
79: data <= 32'Hfffffff2;
80: data <= 32'Hfffffff5;
81: data <= 32'Hfffffff4;
82: data <= 32'Hfffffff2;
83: data <= 32'Hfffffffb;
84: data <= 32'Hfffffff2;
85: data <= 32'Hfffffffd;
86: data <= 32'H00000000;
87: data <= 32'H00000001;
88: data <= 32'H00000006;
89: data <= 32'H00000009;
90: data <= 32'H00000010;
91: data <= 32'H0000000f;
92: data <= 32'H0000000b;
93: data <= 32'H00000011;
94: data <= 32'H0000000f;
95: data <= 32'H0000000b;
96: data <= 32'H0000000f;
97: data <= 32'H00000009;
98: data <= 32'H0000000d;
99: data <= 32'H00000006;
100: data <= 32'H00000003;
101: data <= 32'H00000005;
102: data <= 32'Hffffffff;
103: data <= 32'Hffffffff;
104: data <= 32'Hfffffffa;
105: data <= 32'Hfffffffd;
106: data <= 32'Hfffffffc;
107: data <= 32'Hfffffff9;
108: data <= 32'Hfffffffe;
109: data <= 32'Hfffffffe;
110: data <= 32'Hfffffffd;
111: data <= 32'Hfffffffd;
112: data <= 32'H00000000;
113: data <= 32'Hffffffff;
114: data <= 32'H00000001;
115: data <= 32'H00000006;
116: data <= 32'H00000009;
117: data <= 32'H00000008;
118: data <= 32'H0000000a;
119: data <= 32'H0000000d;
120: data <= 32'H0000000e;
121: data <= 32'H00000015;
122: data <= 32'H00000010;
123: data <= 32'H00000012;
124: data <= 32'H00000013;
125: data <= 32'H0000000f;
126: data <= 32'H0000000f;
127: data <= 32'H00000012;
128: data <= 32'H00000011;
129: data <= 32'Hffffffed;
130: data <= 32'Hfffffff1;
131: data <= 32'Hffffffef;
132: data <= 32'Hffffffea;
133: data <= 32'Hfffffff0;
134: data <= 32'Hfffffff0;
135: data <= 32'Hffffffec;
136: data <= 32'Hfffffff2;
137: data <= 32'Hfffffff1;
138: data <= 32'Hfffffff0;
139: data <= 32'Hfffffff4;
140: data <= 32'Hfffffff4;
141: data <= 32'Hfffffff4;
142: data <= 32'Hfffffff8;
143: data <= 32'Hfffffff5;
144: data <= 32'Hfffffff5;
145: data <= 32'Hfffffff8;
146: data <= 32'Hfffffffb;
147: data <= 32'Hfffffff6;
148: data <= 32'Hfffffff8;
149: data <= 32'Hfffffffb;
150: data <= 32'Hfffffff9;
151: data <= 32'Hfffffffb;
152: data <= 32'Hfffffffc;
153: data <= 32'Hfffffffb;
154: data <= 32'Hfffffffd;
155: data <= 32'Hffffffff;
156: data <= 32'Hfffffff7;
157: data <= 32'Hffffffff;
158: data <= 32'Hfffffffe;
159: data <= 32'Hfffffffa;
160: data <= 32'Hfffffff9;
161: data <= 32'Hfffffffc;
162: data <= 32'Hfffffff7;
163: data <= 32'Hfffffffa;
164: data <= 32'Hfffffff4;
165: data <= 32'Hfffffff8;
166: data <= 32'Hfffffff4;
167: data <= 32'Hfffffff5;
168: data <= 32'Hfffffff4;
169: data <= 32'Hfffffff6;
170: data <= 32'Hfffffff3;
171: data <= 32'Hfffffff4;
172: data <= 32'Hfffffff3;
173: data <= 32'Hfffffff3;
174: data <= 32'Hfffffff4;
175: data <= 32'Hfffffff4;
176: data <= 32'Hfffffffa;
177: data <= 32'Hfffffff9;
178: data <= 32'Hfffffff9;
179: data <= 32'H00000000;
180: data <= 32'Hfffffffd;
181: data <= 32'Hfffffffb;
182: data <= 32'Hffffffff;
183: data <= 32'Hfffffffa;
184: data <= 32'Hfffffff7;
185: data <= 32'Hfffffff5;
186: data <= 32'Hfffffff3;
187: data <= 32'Hffffffee;
188: data <= 32'Hfffffff1;
189: data <= 32'Hffffffef;
190: data <= 32'Hfffffff3;
191: data <= 32'Hfffffff5;
192: data <= 32'Hfffffff6;
193: data <= 32'Hfffffff8;
194: data <= 32'Hfffffff8;
195: data <= 32'Hfffffff8;
196: data <= 32'Hfffffffb;
197: data <= 32'Hfffffffa;
198: data <= 32'Hffffffff;
199: data <= 32'H00000002;
200: data <= 32'Hfffffffd;
201: data <= 32'Hffffffff;
202: data <= 32'H00000002;
203: data <= 32'H00000000;
204: data <= 32'H00000001;
205: data <= 32'H00000001;
206: data <= 32'H00000001;
207: data <= 32'H00000006;
208: data <= 32'H00000004;
209: data <= 32'H00000002;
210: data <= 32'H00000000;
211: data <= 32'H00000002;
212: data <= 32'Hfffffffe;
213: data <= 32'H00000002;
214: data <= 32'Hfffffffe;
215: data <= 32'H00000000;
216: data <= 32'Hfffffffb;
217: data <= 32'H00000005;
218: data <= 32'H00000001;
219: data <= 32'H00000005;
220: data <= 32'H00000004;
221: data <= 32'H00000005;
222: data <= 32'H0000000a;
223: data <= 32'H0000000a;
224: data <= 32'H00000008;
225: data <= 32'H00000009;
226: data <= 32'H00000009;
227: data <= 32'H00000006;
228: data <= 32'H00000007;
229: data <= 32'H0000000a;
230: data <= 32'H0000000c;
231: data <= 32'H0000000a;
232: data <= 32'H0000000f;
233: data <= 32'H0000000c;
234: data <= 32'H00000009;
235: data <= 32'H0000000b;
236: data <= 32'H0000000e;
237: data <= 32'H0000000c;
238: data <= 32'H00000014;
239: data <= 32'H0000000c;
240: data <= 32'H0000000e;
241: data <= 32'H00000009;
242: data <= 32'H00000008;
243: data <= 32'H00000007;
244: data <= 32'H00000009;
245: data <= 32'H00000008;
246: data <= 32'H0000000a;
247: data <= 32'H0000000a;
248: data <= 32'H0000000b;
249: data <= 32'H0000000a;
250: data <= 32'H00000013;
251: data <= 32'H00000013;
252: data <= 32'H00000011;
253: data <= 32'H00000016;
254: data <= 32'H00000011;
255: data <= 32'H00000013;
256: data <= 32'H00000012;
257: data <= 32'Hffffffea;
258: data <= 32'Hffffffec;
259: data <= 32'Hffffffeb;
260: data <= 32'Hffffffee;
261: data <= 32'Hffffffeb;
262: data <= 32'Hfffffff1;
263: data <= 32'Hfffffff0;
264: data <= 32'Hfffffff2;
265: data <= 32'Hfffffff4;
266: data <= 32'Hfffffff7;
267: data <= 32'Hfffffff3;
268: data <= 32'Hfffffffb;
269: data <= 32'Hfffffff7;
270: data <= 32'Hfffffff6;
271: data <= 32'Hfffffff8;
272: data <= 32'Hfffffff9;
273: data <= 32'Hfffffff6;
274: data <= 32'Hfffffffe;
275: data <= 32'Hfffffff9;
276: data <= 32'Hfffffffe;
277: data <= 32'Hfffffffb;
278: data <= 32'Hfffffffe;
279: data <= 32'Hfffffffc;
280: data <= 32'Hfffffffe;
281: data <= 32'Hfffffffd;
282: data <= 32'Hfffffff9;
283: data <= 32'Hfffffffd;
284: data <= 32'Hfffffffc;
285: data <= 32'Hfffffffb;
286: data <= 32'Hfffffffc;
287: data <= 32'Hffffffff;
288: data <= 32'Hfffffff6;
289: data <= 32'Hfffffffd;
290: data <= 32'Hfffffffb;
291: data <= 32'Hfffffff9;
292: data <= 32'Hfffffff7;
293: data <= 32'Hfffffff9;
294: data <= 32'Hfffffff6;
295: data <= 32'Hfffffffc;
296: data <= 32'Hfffffff6;
297: data <= 32'Hfffffff6;
298: data <= 32'Hfffffff3;
299: data <= 32'Hfffffff4;
300: data <= 32'Hfffffff3;
301: data <= 32'Hfffffff5;
302: data <= 32'Hfffffff5;
303: data <= 32'Hfffffffc;
304: data <= 32'Hfffffffc;
305: data <= 32'Hfffffffa;
306: data <= 32'Hfffffffe;
307: data <= 32'Hfffffff9;
308: data <= 32'Hfffffff7;
309: data <= 32'Hfffffff4;
310: data <= 32'Hfffffff2;
311: data <= 32'Hffffffee;
312: data <= 32'Hfffffff0;
313: data <= 32'Hffffffeb;
314: data <= 32'Hffffffee;
315: data <= 32'Hffffffef;
316: data <= 32'Hfffffff1;
317: data <= 32'Hfffffff4;
318: data <= 32'Hfffffff6;
319: data <= 32'Hfffffffc;
320: data <= 32'H00000001;
321: data <= 32'Hffffffff;
322: data <= 32'H00000004;
323: data <= 32'H00000001;
324: data <= 32'H00000002;
325: data <= 32'H0000000f;
326: data <= 32'H0000000e;
327: data <= 32'H00000014;
328: data <= 32'H00000018;
329: data <= 32'H00000011;
330: data <= 32'H00000018;
331: data <= 32'H00000018;
332: data <= 32'H00000012;
333: data <= 32'H00000017;
334: data <= 32'H00000011;
335: data <= 32'H00000011;
336: data <= 32'H0000000b;
337: data <= 32'H0000000a;
338: data <= 32'H00000001;
339: data <= 32'H00000005;
340: data <= 32'Hfffffffd;
341: data <= 32'H00000000;
342: data <= 32'Hfffffff9;
343: data <= 32'H00000000;
344: data <= 32'Hfffffffb;
345: data <= 32'H00000001;
346: data <= 32'Hfffffffc;
347: data <= 32'Hfffffffe;
348: data <= 32'H00000001;
349: data <= 32'H00000005;
350: data <= 32'Hfffffffc;
351: data <= 32'H00000002;
352: data <= 32'Hfffffffd;
353: data <= 32'Hfffffff9;
354: data <= 32'Hfffffffe;
355: data <= 32'Hfffffff6;
356: data <= 32'Hfffffffa;
357: data <= 32'Hfffffffb;
358: data <= 32'Hfffffffe;
359: data <= 32'Hfffffff5;
360: data <= 32'Hffffffff;
361: data <= 32'Hfffffffc;
362: data <= 32'Hfffffffb;
363: data <= 32'Hfffffffa;
364: data <= 32'H00000004;
365: data <= 32'Hffffffff;
366: data <= 32'H0000000f;
367: data <= 32'H00000009;
368: data <= 32'H0000000e;
369: data <= 32'H0000000e;
370: data <= 32'H0000000d;
371: data <= 32'H0000000e;
372: data <= 32'H0000000c;
373: data <= 32'H00000009;
374: data <= 32'H0000000c;
375: data <= 32'H00000008;
376: data <= 32'H00000005;
377: data <= 32'H00000007;
378: data <= 32'H00000009;
379: data <= 32'H00000009;
380: data <= 32'H0000000b;
381: data <= 32'H0000000e;
382: data <= 32'H0000000f;
383: data <= 32'H00000010;
384: data <= 32'H0000000e;
385: data <= 32'Hfffffff3;
386: data <= 32'Hfffffff7;
387: data <= 32'Hfffffff4;
388: data <= 32'Hfffffffa;
389: data <= 32'Hfffffff5;
390: data <= 32'Hfffffffc;
391: data <= 32'Hfffffffb;
392: data <= 32'Hfffffffe;
393: data <= 32'Hfffffffa;
394: data <= 32'H00000000;
395: data <= 32'Hffffffff;
396: data <= 32'Hfffffffe;
397: data <= 32'Hfffffffe;
398: data <= 32'H00000000;
399: data <= 32'Hffffffff;
400: data <= 32'H00000001;
401: data <= 32'H00000001;
402: data <= 32'H00000001;
403: data <= 32'H00000002;
404: data <= 32'H00000003;
405: data <= 32'H00000003;
406: data <= 32'H00000003;
407: data <= 32'H00000005;
408: data <= 32'H00000002;
409: data <= 32'H00000004;
410: data <= 32'Hffffffff;
411: data <= 32'H00000002;
412: data <= 32'H00000001;
413: data <= 32'H00000004;
414: data <= 32'Hfffffffe;
415: data <= 32'H00000007;
416: data <= 32'H00000004;
417: data <= 32'H00000005;
418: data <= 32'H00000002;
419: data <= 32'H00000001;
420: data <= 32'H00000000;
421: data <= 32'H00000004;
422: data <= 32'H00000005;
423: data <= 32'H00000002;
424: data <= 32'H00000001;
425: data <= 32'Hfffffffc;
426: data <= 32'Hfffffffb;
427: data <= 32'Hfffffffb;
428: data <= 32'Hfffffffd;
429: data <= 32'Hfffffff9;
430: data <= 32'H00000000;
431: data <= 32'H00000000;
432: data <= 32'Hfffffffe;
433: data <= 32'Hfffffff9;
434: data <= 32'Hfffffffc;
435: data <= 32'Hfffffff5;
436: data <= 32'Hfffffff1;
437: data <= 32'Hfffffff3;
438: data <= 32'Hfffffff3;
439: data <= 32'Hffffffe8;
440: data <= 32'Hfffffff6;
441: data <= 32'Hfffffff1;
442: data <= 32'Hfffffff6;
443: data <= 32'Hfffffffa;
444: data <= 32'Hfffffffe;
445: data <= 32'Hfffffffd;
446: data <= 32'H00000004;
447: data <= 32'H00000007;
448: data <= 32'H00000009;
449: data <= 32'H0000000c;
450: data <= 32'H0000000c;
451: data <= 32'H0000000b;
452: data <= 32'H0000000e;
453: data <= 32'H0000001b;
454: data <= 32'H00000014;
455: data <= 32'H0000001c;
456: data <= 32'H0000001a;
457: data <= 32'H00000017;
458: data <= 32'H00000015;
459: data <= 32'H0000001a;
460: data <= 32'H00000009;
461: data <= 32'H00000010;
462: data <= 32'H00000009;
463: data <= 32'H00000008;
464: data <= 32'Hfffffffe;
465: data <= 32'H00000003;
466: data <= 32'Hffffffff;
467: data <= 32'Hfffffffb;
468: data <= 32'Hfffffff7;
469: data <= 32'Hfffffffd;
470: data <= 32'Hfffffff9;
471: data <= 32'H00000003;
472: data <= 32'Hfffffffc;
473: data <= 32'H00000004;
474: data <= 32'H00000001;
475: data <= 32'H00000004;
476: data <= 32'H0000000a;
477: data <= 32'H0000000c;
478: data <= 32'H00000004;
479: data <= 32'H00000001;
480: data <= 32'H00000000;
481: data <= 32'Hfffffffa;
482: data <= 32'H00000001;
483: data <= 32'Hfffffffa;
484: data <= 32'H00000001;
485: data <= 32'Hfffffffb;
486: data <= 32'H00000001;
487: data <= 32'Hfffffff6;
488: data <= 32'Hfffffffd;
489: data <= 32'Hfffffff8;
490: data <= 32'Hfffffff3;
491: data <= 32'Hfffffff1;
492: data <= 32'Hfffffff2;
493: data <= 32'Hffffffeb;
494: data <= 32'Hfffffff9;
495: data <= 32'Hfffffff7;
496: data <= 32'Hfffffffc;
497: data <= 32'H00000002;
498: data <= 32'H00000005;
499: data <= 32'H0000000e;
500: data <= 32'H0000000a;
501: data <= 32'H00000012;
502: data <= 32'H00000014;
503: data <= 32'H0000000d;
504: data <= 32'H00000010;
505: data <= 32'H00000011;
506: data <= 32'H0000000b;
507: data <= 32'H0000000e;
508: data <= 32'H0000000d;
509: data <= 32'H0000000f;
510: data <= 32'H0000000e;
511: data <= 32'H00000016;
512: data <= 32'H00000010;
513: data <= 32'Hfffffffe;
514: data <= 32'Hffffffff;
515: data <= 32'Hfffffffe;
516: data <= 32'H00000002;
517: data <= 32'Hfffffffd;
518: data <= 32'H00000002;
519: data <= 32'H00000002;
520: data <= 32'H00000004;
521: data <= 32'H00000002;
522: data <= 32'H00000006;
523: data <= 32'H00000004;
524: data <= 32'H00000005;
525: data <= 32'H00000004;
526: data <= 32'H0000000a;
527: data <= 32'H00000007;
528: data <= 32'H00000009;
529: data <= 32'H0000000b;
530: data <= 32'H00000007;
531: data <= 32'H00000007;
532: data <= 32'H00000006;
533: data <= 32'H0000000a;
534: data <= 32'H00000006;
535: data <= 32'H0000000b;
536: data <= 32'H00000005;
537: data <= 32'H0000000c;
538: data <= 32'H00000007;
539: data <= 32'H0000000b;
540: data <= 32'H00000007;
541: data <= 32'H0000000d;
542: data <= 32'H00000008;
543: data <= 32'H0000000e;
544: data <= 32'H0000000e;
545: data <= 32'H0000000e;
546: data <= 32'H0000000a;
547: data <= 32'H0000000b;
548: data <= 32'H00000009;
549: data <= 32'H0000000d;
550: data <= 32'H0000000e;
551: data <= 32'H00000008;
552: data <= 32'H00000006;
553: data <= 32'H00000004;
554: data <= 32'H00000002;
555: data <= 32'H00000001;
556: data <= 32'H00000004;
557: data <= 32'Hfffffffe;
558: data <= 32'H00000008;
559: data <= 32'H00000002;
560: data <= 32'Hfffffffc;
561: data <= 32'Hfffffff7;
562: data <= 32'Hfffffffb;
563: data <= 32'Hfffffff0;
564: data <= 32'Hfffffff4;
565: data <= 32'Hfffffff3;
566: data <= 32'Hfffffff9;
567: data <= 32'Hfffffff5;
568: data <= 32'Hffffffff;
569: data <= 32'H00000000;
570: data <= 32'H00000003;
571: data <= 32'H00000003;
572: data <= 32'H00000009;
573: data <= 32'H00000006;
574: data <= 32'H00000006;
575: data <= 32'H0000000c;
576: data <= 32'H00000009;
577: data <= 32'H0000000e;
578: data <= 32'H00000011;
579: data <= 32'H0000000f;
580: data <= 32'H00000011;
581: data <= 32'H00000018;
582: data <= 32'H00000012;
583: data <= 32'H00000015;
584: data <= 32'H00000012;
585: data <= 32'H0000000f;
586: data <= 32'H0000000e;
587: data <= 32'H0000000f;
588: data <= 32'H00000000;
589: data <= 32'H00000006;
590: data <= 32'H00000001;
591: data <= 32'H00000003;
592: data <= 32'Hfffffff9;
593: data <= 32'Hfffffffe;
594: data <= 32'Hfffffffa;
595: data <= 32'Hfffffff7;
596: data <= 32'Hfffffff5;
597: data <= 32'Hfffffffb;
598: data <= 32'Hfffffffa;
599: data <= 32'Hfffffffd;
600: data <= 32'Hfffffffd;
601: data <= 32'Hfffffffe;
602: data <= 32'H00000000;
603: data <= 32'H00000003;
604: data <= 32'H00000007;
605: data <= 32'H00000000;
606: data <= 32'Hfffffff4;
607: data <= 32'Hfffffff1;
608: data <= 32'Hffffffec;
609: data <= 32'Hffffffe5;
610: data <= 32'Hfffffff1;
611: data <= 32'Hffffffec;
612: data <= 32'Hfffffff7;
613: data <= 32'Hfffffff5;
614: data <= 32'H00000000;
615: data <= 32'H00000005;
616: data <= 32'H00000006;
617: data <= 32'H00000005;
618: data <= 32'H00000006;
619: data <= 32'Hffffffff;
620: data <= 32'Hfffffff8;
621: data <= 32'Hfffffff4;
622: data <= 32'Hfffffff6;
623: data <= 32'Hffffffee;
624: data <= 32'Hfffffff0;
625: data <= 32'Hfffffff4;
626: data <= 32'Hfffffff0;
627: data <= 32'Hfffffffe;
628: data <= 32'Hffffffff;
629: data <= 32'H00000006;
630: data <= 32'H0000000c;
631: data <= 32'H0000000d;
632: data <= 32'H0000000d;
633: data <= 32'H00000017;
634: data <= 32'H00000010;
635: data <= 32'H00000015;
636: data <= 32'H00000014;
637: data <= 32'H00000014;
638: data <= 32'H00000012;
639: data <= 32'H0000001b;
640: data <= 32'H00000018;
641: data <= 32'Hfffffff6;
642: data <= 32'Hfffffffa;
643: data <= 32'Hfffffff8;
644: data <= 32'Hfffffffa;
645: data <= 32'Hfffffff8;
646: data <= 32'Hfffffffa;
647: data <= 32'Hfffffffe;
648: data <= 32'Hfffffffd;
649: data <= 32'Hffffffff;
650: data <= 32'H00000003;
651: data <= 32'Hfffffffd;
652: data <= 32'H00000005;
653: data <= 32'H00000003;
654: data <= 32'H00000003;
655: data <= 32'H00000006;
656: data <= 32'H00000006;
657: data <= 32'H00000006;
658: data <= 32'H00000005;
659: data <= 32'H00000005;
660: data <= 32'Hffffffff;
661: data <= 32'H00000005;
662: data <= 32'H00000004;
663: data <= 32'H00000000;
664: data <= 32'H00000001;
665: data <= 32'H00000006;
666: data <= 32'H00000004;
667: data <= 32'H00000006;
668: data <= 32'H00000006;
669: data <= 32'H00000005;
670: data <= 32'H00000007;
671: data <= 32'H00000007;
672: data <= 32'H00000004;
673: data <= 32'H00000006;
674: data <= 32'H00000002;
675: data <= 32'H00000004;
676: data <= 32'H00000002;
677: data <= 32'H00000005;
678: data <= 32'H00000003;
679: data <= 32'H00000000;
680: data <= 32'Hfffffffd;
681: data <= 32'Hfffffffd;
682: data <= 32'Hfffffffa;
683: data <= 32'Hfffffff8;
684: data <= 32'Hfffffff8;
685: data <= 32'Hfffffff3;
686: data <= 32'Hfffffff4;
687: data <= 32'Hfffffff7;
688: data <= 32'Hfffffff6;
689: data <= 32'Hfffffff1;
690: data <= 32'Hfffffff9;
691: data <= 32'Hfffffff8;
692: data <= 32'Hfffffff6;
693: data <= 32'H00000000;
694: data <= 32'H00000001;
695: data <= 32'Hfffffffd;
696: data <= 32'H00000002;
697: data <= 32'Hffffffff;
698: data <= 32'Hfffffffb;
699: data <= 32'Hfffffffb;
700: data <= 32'H00000001;
701: data <= 32'Hfffffffb;
702: data <= 32'Hfffffffe;
703: data <= 32'H00000003;
704: data <= 32'Hfffffffe;
705: data <= 32'H00000000;
706: data <= 32'H00000001;
707: data <= 32'Hfffffffb;
708: data <= 32'Hfffffffc;
709: data <= 32'Hfffffffd;
710: data <= 32'Hfffffffb;
711: data <= 32'H00000000;
712: data <= 32'H00000001;
713: data <= 32'H00000004;
714: data <= 32'H0000000b;
715: data <= 32'H00000007;
716: data <= 32'H00000002;
717: data <= 32'H00000008;
718: data <= 32'H00000003;
719: data <= 32'H00000004;
720: data <= 32'H00000000;
721: data <= 32'H00000000;
722: data <= 32'Hfffffffe;
723: data <= 32'H00000001;
724: data <= 32'H00000002;
725: data <= 32'H00000007;
726: data <= 32'H00000007;
727: data <= 32'H00000008;
728: data <= 32'H00000006;
729: data <= 32'H00000006;
730: data <= 32'H00000001;
731: data <= 32'Hffffffff;
732: data <= 32'Hfffffffc;
733: data <= 32'Hffffffed;
734: data <= 32'Hffffffe3;
735: data <= 32'Hffffffe0;
736: data <= 32'Hffffffd8;
737: data <= 32'Hffffffcd;
738: data <= 32'Hffffffcf;
739: data <= 32'Hffffffcb;
740: data <= 32'Hffffffce;
741: data <= 32'Hffffffd0;
742: data <= 32'Hffffffe5;
743: data <= 32'Hfffffff1;
744: data <= 32'Hfffffff5;
745: data <= 32'H00000002;
746: data <= 32'H00000008;
747: data <= 32'H00000005;
748: data <= 32'H00000000;
749: data <= 32'H00000003;
750: data <= 32'Hffffffff;
751: data <= 32'Hfffffff3;
752: data <= 32'Hfffffff4;
753: data <= 32'Hfffffff3;
754: data <= 32'Hffffffe6;
755: data <= 32'Hffffffee;
756: data <= 32'Hfffffff0;
757: data <= 32'Hffffffeb;
758: data <= 32'Hfffffff2;
759: data <= 32'Hfffffff5;
760: data <= 32'Hfffffff9;
761: data <= 32'H00000004;
762: data <= 32'H00000005;
763: data <= 32'H00000009;
764: data <= 32'H0000000f;
765: data <= 32'H0000000c;
766: data <= 32'H0000000c;
767: data <= 32'H00000012;
768: data <= 32'H00000010;
769: data <= 32'H00000000;
770: data <= 32'H00000001;
771: data <= 32'H00000004;
772: data <= 32'Hfffffffe;
773: data <= 32'H00000006;
774: data <= 32'H00000003;
775: data <= 32'H00000005;
776: data <= 32'H0000000a;
777: data <= 32'H00000009;
778: data <= 32'H00000008;
779: data <= 32'H00000010;
780: data <= 32'H0000000c;
781: data <= 32'H00000009;
782: data <= 32'H00000010;
783: data <= 32'H0000000d;
784: data <= 32'H0000000a;
785: data <= 32'H00000011;
786: data <= 32'H0000000e;
787: data <= 32'H0000000b;
788: data <= 32'H0000000e;
789: data <= 32'H0000000b;
790: data <= 32'H0000000b;
791: data <= 32'H0000000b;
792: data <= 32'H0000000d;
793: data <= 32'H0000000b;
794: data <= 32'H0000000f;
795: data <= 32'H0000000c;
796: data <= 32'H00000010;
797: data <= 32'H0000000d;
798: data <= 32'H00000010;
799: data <= 32'H0000000b;
800: data <= 32'H00000010;
801: data <= 32'H00000010;
802: data <= 32'H00000011;
803: data <= 32'H00000014;
804: data <= 32'H00000013;
805: data <= 32'H00000014;
806: data <= 32'H00000015;
807: data <= 32'H0000000c;
808: data <= 32'H00000008;
809: data <= 32'H00000008;
810: data <= 32'H00000001;
811: data <= 32'H00000003;
812: data <= 32'Hfffffffe;
813: data <= 32'Hfffffffc;
814: data <= 32'H00000001;
815: data <= 32'H00000007;
816: data <= 32'H00000004;
817: data <= 32'H00000009;
818: data <= 32'H00000006;
819: data <= 32'H00000009;
820: data <= 32'H00000006;
821: data <= 32'H00000009;
822: data <= 32'H0000000a;
823: data <= 32'H00000008;
824: data <= 32'H00000008;
825: data <= 32'H0000000d;
826: data <= 32'H00000004;
827: data <= 32'H00000009;
828: data <= 32'H00000008;
829: data <= 32'Hffffffff;
830: data <= 32'Hfffffffc;
831: data <= 32'Hfffffffc;
832: data <= 32'Hfffffff3;
833: data <= 32'Hfffffff1;
834: data <= 32'Hfffffff0;
835: data <= 32'Hffffffee;
836: data <= 32'Hffffffef;
837: data <= 32'Hfffffff7;
838: data <= 32'Hfffffff7;
839: data <= 32'Hfffffffc;
840: data <= 32'Hffffffff;
841: data <= 32'H00000000;
842: data <= 32'H00000006;
843: data <= 32'Hfffffffb;
844: data <= 32'Hfffffffb;
845: data <= 32'Hfffffff3;
846: data <= 32'Hfffffff4;
847: data <= 32'Hfffffff4;
848: data <= 32'Hfffffff5;
849: data <= 32'Hfffffff4;
850: data <= 32'Hfffffff6;
851: data <= 32'Hfffffffa;
852: data <= 32'H00000001;
853: data <= 32'H0000000a;
854: data <= 32'H0000000f;
855: data <= 32'H00000015;
856: data <= 32'H00000017;
857: data <= 32'H00000017;
858: data <= 32'H00000016;
859: data <= 32'H00000012;
860: data <= 32'H0000000c;
861: data <= 32'H00000007;
862: data <= 32'H00000002;
863: data <= 32'H00000003;
864: data <= 32'Hfffffffb;
865: data <= 32'Hffffffee;
866: data <= 32'Hffffffe4;
867: data <= 32'Hffffffd8;
868: data <= 32'Hffffffd3;
869: data <= 32'Hffffffcf;
870: data <= 32'Hffffffdc;
871: data <= 32'Hfffffff1;
872: data <= 32'Hfffffff2;
873: data <= 32'Hfffffffa;
874: data <= 32'Hfffffffc;
875: data <= 32'Hfffffffd;
876: data <= 32'Hfffffffa;
877: data <= 32'H00000004;
878: data <= 32'H00000002;
879: data <= 32'H00000002;
880: data <= 32'H00000008;
881: data <= 32'H00000005;
882: data <= 32'Hffffffff;
883: data <= 32'Hffffffff;
884: data <= 32'Hfffffffd;
885: data <= 32'Hfffffff6;
886: data <= 32'Hfffffff3;
887: data <= 32'Hfffffff4;
888: data <= 32'Hfffffff8;
889: data <= 32'Hfffffff6;
890: data <= 32'Hfffffffe;
891: data <= 32'H00000002;
892: data <= 32'H00000007;
893: data <= 32'H0000000d;
894: data <= 32'H00000012;
895: data <= 32'H00000010;
896: data <= 32'H00000012;
897: data <= 32'H00000005;
898: data <= 32'H00000005;
899: data <= 32'H0000000a;
900: data <= 32'H00000007;
901: data <= 32'H0000000a;
902: data <= 32'H00000006;
903: data <= 32'H0000000e;
904: data <= 32'H00000008;
905: data <= 32'H00000011;
906: data <= 32'H00000013;
907: data <= 32'H00000013;
908: data <= 32'H00000018;
909: data <= 32'H00000016;
910: data <= 32'H0000000f;
911: data <= 32'H00000016;
912: data <= 32'H00000015;
913: data <= 32'H00000013;
914: data <= 32'H00000012;
915: data <= 32'H00000012;
916: data <= 32'H00000013;
917: data <= 32'H00000012;
918: data <= 32'H00000016;
919: data <= 32'H00000011;
920: data <= 32'H00000013;
921: data <= 32'H00000012;
922: data <= 32'H0000000e;
923: data <= 32'H0000000c;
924: data <= 32'H00000017;
925: data <= 32'H0000000c;
926: data <= 32'H00000017;
927: data <= 32'H00000014;
928: data <= 32'H00000014;
929: data <= 32'H00000017;
930: data <= 32'H00000016;
931: data <= 32'H00000013;
932: data <= 32'H00000018;
933: data <= 32'H00000013;
934: data <= 32'H00000016;
935: data <= 32'H0000000b;
936: data <= 32'H00000006;
937: data <= 32'H00000003;
938: data <= 32'Hfffffffe;
939: data <= 32'Hfffffff9;
940: data <= 32'Hfffffffa;
941: data <= 32'Hfffffffc;
942: data <= 32'Hfffffffa;
943: data <= 32'H00000006;
944: data <= 32'Hfffffffe;
945: data <= 32'H00000002;
946: data <= 32'H00000002;
947: data <= 32'H00000001;
948: data <= 32'Hfffffffd;
949: data <= 32'H00000005;
950: data <= 32'Hfffffffb;
951: data <= 32'Hfffffff9;
952: data <= 32'Hffffffff;
953: data <= 32'Hfffffff6;
954: data <= 32'Hffffffeb;
955: data <= 32'Hffffffef;
956: data <= 32'Hffffffec;
957: data <= 32'Hffffffe7;
958: data <= 32'Hffffffe4;
959: data <= 32'Hffffffea;
960: data <= 32'Hffffffe9;
961: data <= 32'Hffffffe7;
962: data <= 32'Hffffffed;
963: data <= 32'Hfffffff5;
964: data <= 32'Hfffffff7;
965: data <= 32'Hfffffffd;
966: data <= 32'H00000000;
967: data <= 32'Hffffffff;
968: data <= 32'H00000006;
969: data <= 32'Hfffffffe;
970: data <= 32'H00000006;
971: data <= 32'Hfffffffa;
972: data <= 32'H00000000;
973: data <= 32'Hfffffffd;
974: data <= 32'Hfffffffb;
975: data <= 32'Hfffffffd;
976: data <= 32'H00000005;
977: data <= 32'Hffffffff;
978: data <= 32'H00000004;
979: data <= 32'H00000007;
980: data <= 32'H0000000e;
981: data <= 32'H0000000b;
982: data <= 32'H00000011;
983: data <= 32'H00000011;
984: data <= 32'H00000013;
985: data <= 32'H00000010;
986: data <= 32'H0000000c;
987: data <= 32'H0000000c;
988: data <= 32'H00000006;
989: data <= 32'H00000004;
990: data <= 32'H00000005;
991: data <= 32'H00000008;
992: data <= 32'H00000008;
993: data <= 32'Hfffffffc;
994: data <= 32'Hfffffff6;
995: data <= 32'Hffffffee;
996: data <= 32'Hffffffe4;
997: data <= 32'Hffffffe2;
998: data <= 32'Hffffffef;
999: data <= 32'Hfffffffc;
1000: data <= 32'Hfffffffc;
1001: data <= 32'Hfffffffe;
1002: data <= 32'Hfffffffb;
1003: data <= 32'Hfffffffc;
1004: data <= 32'Hfffffff0;
1005: data <= 32'Hfffffff9;
1006: data <= 32'Hfffffff1;
1007: data <= 32'Hfffffff5;
1008: data <= 32'Hfffffff5;
1009: data <= 32'Hfffffffd;
1010: data <= 32'Hfffffff5;
1011: data <= 32'Hfffffff9;
1012: data <= 32'Hfffffffc;
1013: data <= 32'Hfffffff5;
1014: data <= 32'Hfffffffb;
1015: data <= 32'Hfffffff9;
1016: data <= 32'Hfffffffb;
1017: data <= 32'Hfffffffb;
1018: data <= 32'Hfffffff7;
1019: data <= 32'Hfffffff9;
1020: data <= 32'Hfffffffe;
1021: data <= 32'Hfffffffa;
1022: data <= 32'H0000000a;
1023: data <= 32'H00000006;
1024: data <= 32'H0000000f;
1025: data <= 32'Hfffffffc;
1026: data <= 32'Hfffffffc;
1027: data <= 32'H00000000;
1028: data <= 32'Hfffffffa;
1029: data <= 32'H00000002;
1030: data <= 32'Hfffffffe;
1031: data <= 32'H00000000;
1032: data <= 32'H00000003;
1033: data <= 32'H00000002;
1034: data <= 32'H00000006;
1035: data <= 32'H00000008;
1036: data <= 32'H00000009;
1037: data <= 32'H00000008;
1038: data <= 32'H0000000b;
1039: data <= 32'H0000000a;
1040: data <= 32'H0000000a;
1041: data <= 32'H0000000c;
1042: data <= 32'H00000005;
1043: data <= 32'H00000006;
1044: data <= 32'H00000006;
1045: data <= 32'H00000009;
1046: data <= 32'H00000006;
1047: data <= 32'H00000007;
1048: data <= 32'H00000007;
1049: data <= 32'H00000005;
1050: data <= 32'H00000006;
1051: data <= 32'H00000007;
1052: data <= 32'H00000009;
1053: data <= 32'H00000009;
1054: data <= 32'H0000000b;
1055: data <= 32'H0000000c;
1056: data <= 32'H00000010;
1057: data <= 32'H0000000f;
1058: data <= 32'H00000010;
1059: data <= 32'H00000013;
1060: data <= 32'H0000000c;
1061: data <= 32'H0000000b;
1062: data <= 32'H00000008;
1063: data <= 32'Hfffffff8;
1064: data <= 32'Hfffffffa;
1065: data <= 32'Hfffffff6;
1066: data <= 32'Hffffffef;
1067: data <= 32'Hfffffff4;
1068: data <= 32'Hfffffff5;
1069: data <= 32'Hffffffed;
1070: data <= 32'Hffffffee;
1071: data <= 32'Hfffffff3;
1072: data <= 32'Hffffffea;
1073: data <= 32'Hffffffef;
1074: data <= 32'Hffffffee;
1075: data <= 32'Hffffffef;
1076: data <= 32'Hffffffea;
1077: data <= 32'Hffffffef;
1078: data <= 32'Hffffffe9;
1079: data <= 32'Hffffffe1;
1080: data <= 32'Hffffffe6;
1081: data <= 32'Hffffffe5;
1082: data <= 32'Hffffffd9;
1083: data <= 32'Hffffffde;
1084: data <= 32'Hffffffde;
1085: data <= 32'Hffffffdd;
1086: data <= 32'Hffffffe6;
1087: data <= 32'Hffffffef;
1088: data <= 32'Hfffffff4;
1089: data <= 32'H00000000;
1090: data <= 32'H00000003;
1091: data <= 32'H00000004;
1092: data <= 32'H0000000d;
1093: data <= 32'H0000000a;
1094: data <= 32'H0000000d;
1095: data <= 32'H0000000d;
1096: data <= 32'H00000011;
1097: data <= 32'H00000016;
1098: data <= 32'H0000001a;
1099: data <= 32'H00000012;
1100: data <= 32'H00000014;
1101: data <= 32'H0000000b;
1102: data <= 32'H00000001;
1103: data <= 32'Hfffffffa;
1104: data <= 32'Hfffffffa;
1105: data <= 32'Hffffffee;
1106: data <= 32'Hffffffe9;
1107: data <= 32'Hffffffe6;
1108: data <= 32'Hffffffe7;
1109: data <= 32'Hffffffe4;
1110: data <= 32'Hffffffe5;
1111: data <= 32'Hffffffe8;
1112: data <= 32'Hffffffeb;
1113: data <= 32'Hffffffee;
1114: data <= 32'Hffffffed;
1115: data <= 32'Hfffffff3;
1116: data <= 32'Hfffffff1;
1117: data <= 32'Hfffffff2;
1118: data <= 32'Hfffffff5;
1119: data <= 32'Hfffffff9;
1120: data <= 32'Hfffffff5;
1121: data <= 32'Hfffffff3;
1122: data <= 32'Hfffffff4;
1123: data <= 32'Hfffffff4;
1124: data <= 32'Hfffffff1;
1125: data <= 32'Hfffffff1;
1126: data <= 32'Hfffffff8;
1127: data <= 32'Hffffffff;
1128: data <= 32'H00000000;
1129: data <= 32'H00000003;
1130: data <= 32'H00000000;
1131: data <= 32'Hfffffffe;
1132: data <= 32'Hfffffff3;
1133: data <= 32'Hfffffff1;
1134: data <= 32'Hffffffeb;
1135: data <= 32'Hffffffec;
1136: data <= 32'Hffffffe7;
1137: data <= 32'Hffffffed;
1138: data <= 32'Hffffffe8;
1139: data <= 32'Hffffffe3;
1140: data <= 32'Hffffffe3;
1141: data <= 32'Hffffffe7;
1142: data <= 32'Hffffffe2;
1143: data <= 32'Hffffffe7;
1144: data <= 32'Hffffffee;
1145: data <= 32'Hffffffed;
1146: data <= 32'Hfffffff0;
1147: data <= 32'Hfffffff4;
1148: data <= 32'Hfffffffb;
1149: data <= 32'Hfffffff1;
1150: data <= 32'Hfffffff8;
1151: data <= 32'Hfffffff8;
1152: data <= 32'Hfffffffd;
1153: data <= 32'Hfffffff8;
1154: data <= 32'Hfffffff4;
1155: data <= 32'Hfffffff6;
1156: data <= 32'Hfffffff4;
1157: data <= 32'Hfffffff4;
1158: data <= 32'Hfffffff6;
1159: data <= 32'Hfffffff5;
1160: data <= 32'Hfffffffb;
1161: data <= 32'Hfffffff8;
1162: data <= 32'H00000000;
1163: data <= 32'Hfffffffb;
1164: data <= 32'H00000001;
1165: data <= 32'Hfffffffb;
1166: data <= 32'H00000002;
1167: data <= 32'H00000002;
1168: data <= 32'H00000000;
1169: data <= 32'Hffffffff;
1170: data <= 32'H00000000;
1171: data <= 32'H00000001;
1172: data <= 32'Hfffffffa;
1173: data <= 32'H00000001;
1174: data <= 32'Hfffffffe;
1175: data <= 32'Hfffffffa;
1176: data <= 32'Hfffffffe;
1177: data <= 32'Hfffffffc;
1178: data <= 32'Hfffffffa;
1179: data <= 32'Hffffffff;
1180: data <= 32'H00000000;
1181: data <= 32'H00000002;
1182: data <= 32'H00000004;
1183: data <= 32'H00000006;
1184: data <= 32'H00000004;
1185: data <= 32'H00000006;
1186: data <= 32'H00000002;
1187: data <= 32'H00000004;
1188: data <= 32'H00000000;
1189: data <= 32'Hfffffffc;
1190: data <= 32'Hfffffff8;
1191: data <= 32'Hfffffff6;
1192: data <= 32'Hfffffff0;
1193: data <= 32'Hffffffef;
1194: data <= 32'Hffffffe7;
1195: data <= 32'Hffffffe1;
1196: data <= 32'Hffffffe1;
1197: data <= 32'Hffffffdb;
1198: data <= 32'Hffffffe7;
1199: data <= 32'Hfffffff6;
1200: data <= 32'Hffffffee;
1201: data <= 32'Hfffffff4;
1202: data <= 32'Hfffffff6;
1203: data <= 32'Hffffffe8;
1204: data <= 32'Hffffffe7;
1205: data <= 32'Hffffffe5;
1206: data <= 32'Hffffffdd;
1207: data <= 32'Hffffffdc;
1208: data <= 32'Hffffffe0;
1209: data <= 32'Hffffffe0;
1210: data <= 32'Hffffffe4;
1211: data <= 32'Hffffffe7;
1212: data <= 32'Hffffffed;
1213: data <= 32'Hfffffff7;
1214: data <= 32'Hffffffff;
1215: data <= 32'H0000000a;
1216: data <= 32'H00000011;
1217: data <= 32'H00000012;
1218: data <= 32'H00000013;
1219: data <= 32'H00000010;
1220: data <= 32'H00000018;
1221: data <= 32'H0000001d;
1222: data <= 32'H00000017;
1223: data <= 32'H00000018;
1224: data <= 32'H00000018;
1225: data <= 32'H00000010;
1226: data <= 32'H00000008;
1227: data <= 32'H00000003;
1228: data <= 32'Hfffffffb;
1229: data <= 32'Hfffffff7;
1230: data <= 32'Hfffffff2;
1231: data <= 32'Hfffffff2;
1232: data <= 32'Hfffffff3;
1233: data <= 32'Hfffffff1;
1234: data <= 32'Hffffffec;
1235: data <= 32'Hffffffef;
1236: data <= 32'Hffffffec;
1237: data <= 32'Hffffffee;
1238: data <= 32'Hffffffe9;
1239: data <= 32'Hffffffef;
1240: data <= 32'Hffffffec;
1241: data <= 32'Hffffffee;
1242: data <= 32'Hffffffed;
1243: data <= 32'Hfffffff0;
1244: data <= 32'Hfffffff0;
1245: data <= 32'Hfffffff5;
1246: data <= 32'Hfffffff8;
1247: data <= 32'Hfffffffa;
1248: data <= 32'Hffffffff;
1249: data <= 32'Hfffffffd;
1250: data <= 32'H00000002;
1251: data <= 32'Hfffffffe;
1252: data <= 32'Hfffffffd;
1253: data <= 32'H00000002;
1254: data <= 32'H00000000;
1255: data <= 32'Hfffffffd;
1256: data <= 32'H00000004;
1257: data <= 32'H00000000;
1258: data <= 32'H00000009;
1259: data <= 32'H00000007;
1260: data <= 32'H00000004;
1261: data <= 32'Hfffffffd;
1262: data <= 32'Hfffffff5;
1263: data <= 32'Hfffffff2;
1264: data <= 32'Hffffffed;
1265: data <= 32'Hffffffec;
1266: data <= 32'Hffffffea;
1267: data <= 32'Hffffffe4;
1268: data <= 32'Hffffffe5;
1269: data <= 32'Hffffffe7;
1270: data <= 32'Hffffffe6;
1271: data <= 32'Hffffffe8;
1272: data <= 32'Hffffffea;
1273: data <= 32'Hffffffec;
1274: data <= 32'Hffffffea;
1275: data <= 32'Hffffffef;
1276: data <= 32'Hfffffff7;
1277: data <= 32'Hfffffff5;
1278: data <= 32'Hfffffff9;
1279: data <= 32'H00000000;
1280: data <= 32'H00000000;
1281: data <= 32'H00000003;
1282: data <= 32'H00000002;
1283: data <= 32'Hffffffff;
1284: data <= 32'H00000002;
1285: data <= 32'Hfffffffd;
1286: data <= 32'H00000003;
1287: data <= 32'Hfffffffe;
1288: data <= 32'H00000006;
1289: data <= 32'H00000001;
1290: data <= 32'H00000009;
1291: data <= 32'H00000005;
1292: data <= 32'H00000009;
1293: data <= 32'H00000005;
1294: data <= 32'H0000000a;
1295: data <= 32'H00000006;
1296: data <= 32'H00000009;
1297: data <= 32'H00000007;
1298: data <= 32'H00000008;
1299: data <= 32'H00000008;
1300: data <= 32'H00000003;
1301: data <= 32'H00000008;
1302: data <= 32'H00000004;
1303: data <= 32'H00000000;
1304: data <= 32'H00000001;
1305: data <= 32'H00000002;
1306: data <= 32'Hfffffffe;
1307: data <= 32'H00000004;
1308: data <= 32'H00000007;
1309: data <= 32'H0000000c;
1310: data <= 32'H00000007;
1311: data <= 32'H0000000c;
1312: data <= 32'H00000002;
1313: data <= 32'H00000003;
1314: data <= 32'H00000003;
1315: data <= 32'H00000007;
1316: data <= 32'H00000002;
1317: data <= 32'H00000004;
1318: data <= 32'Hfffffffe;
1319: data <= 32'Hfffffff3;
1320: data <= 32'Hfffffff1;
1321: data <= 32'Hffffffef;
1322: data <= 32'Hffffffe6;
1323: data <= 32'Hffffffec;
1324: data <= 32'Hfffffff6;
1325: data <= 32'Hfffffffc;
1326: data <= 32'H00000006;
1327: data <= 32'H00000009;
1328: data <= 32'Hffffffff;
1329: data <= 32'Hfffffffe;
1330: data <= 32'Hfffffff8;
1331: data <= 32'Hffffffea;
1332: data <= 32'Hffffffea;
1333: data <= 32'Hffffffeb;
1334: data <= 32'Hffffffee;
1335: data <= 32'Hffffffee;
1336: data <= 32'Hfffffffc;
1337: data <= 32'Hfffffffe;
1338: data <= 32'H00000002;
1339: data <= 32'H00000003;
1340: data <= 32'H0000000c;
1341: data <= 32'H0000000b;
1342: data <= 32'H00000012;
1343: data <= 32'H00000015;
1344: data <= 32'H00000013;
1345: data <= 32'H00000012;
1346: data <= 32'H0000000b;
1347: data <= 32'H00000009;
1348: data <= 32'H0000000c;
1349: data <= 32'H00000009;
1350: data <= 32'H00000003;
1351: data <= 32'H00000009;
1352: data <= 32'H00000003;
1353: data <= 32'H00000003;
1354: data <= 32'Hfffffffb;
1355: data <= 32'Hfffffffd;
1356: data <= 32'Hfffffffa;
1357: data <= 32'Hffffffff;
1358: data <= 32'Hfffffffd;
1359: data <= 32'Hffffffff;
1360: data <= 32'Hfffffffc;
1361: data <= 32'Hfffffffe;
1362: data <= 32'Hfffffffa;
1363: data <= 32'Hfffffffe;
1364: data <= 32'Hfffffff8;
1365: data <= 32'Hfffffffb;
1366: data <= 32'Hfffffff7;
1367: data <= 32'Hfffffff6;
1368: data <= 32'Hfffffff1;
1369: data <= 32'Hfffffff5;
1370: data <= 32'Hfffffff0;
1371: data <= 32'Hfffffff2;
1372: data <= 32'Hffffffec;
1373: data <= 32'Hffffffea;
1374: data <= 32'Hffffffec;
1375: data <= 32'Hffffffec;
1376: data <= 32'Hfffffff2;
1377: data <= 32'Hfffffff5;
1378: data <= 32'Hfffffffa;
1379: data <= 32'Hfffffff9;
1380: data <= 32'Hfffffffb;
1381: data <= 32'Hfffffffa;
1382: data <= 32'Hfffffffe;
1383: data <= 32'Hfffffff9;
1384: data <= 32'H00000000;
1385: data <= 32'Hfffffffe;
1386: data <= 32'H00000001;
1387: data <= 32'H00000002;
1388: data <= 32'H00000006;
1389: data <= 32'Hfffffffa;
1390: data <= 32'Hfffffffa;
1391: data <= 32'Hfffffff9;
1392: data <= 32'Hfffffff5;
1393: data <= 32'Hfffffff3;
1394: data <= 32'Hfffffff7;
1395: data <= 32'Hffffffea;
1396: data <= 32'Hffffffe9;
1397: data <= 32'Hfffffff1;
1398: data <= 32'Hffffffef;
1399: data <= 32'Hfffffff4;
1400: data <= 32'Hfffffffd;
1401: data <= 32'Hffffffff;
1402: data <= 32'Hfffffffd;
1403: data <= 32'H00000002;
1404: data <= 32'H00000001;
1405: data <= 32'H00000002;
1406: data <= 32'H00000004;
1407: data <= 32'H0000000c;
1408: data <= 32'H0000000c;
1409: data <= 32'H00000006;
1410: data <= 32'H00000001;
1411: data <= 32'Hfffffffe;
1412: data <= 32'H00000003;
1413: data <= 32'Hffffffff;
1414: data <= 32'H00000000;
1415: data <= 32'H00000000;
1416: data <= 32'H00000003;
1417: data <= 32'Hffffffff;
1418: data <= 32'H00000006;
1419: data <= 32'H00000006;
1420: data <= 32'H00000005;
1421: data <= 32'H00000005;
1422: data <= 32'H00000008;
1423: data <= 32'H00000002;
1424: data <= 32'H00000008;
1425: data <= 32'H00000009;
1426: data <= 32'H00000005;
1427: data <= 32'H00000002;
1428: data <= 32'H00000001;
1429: data <= 32'Hffffffff;
1430: data <= 32'H00000001;
1431: data <= 32'Hffffffff;
1432: data <= 32'Hfffffffd;
1433: data <= 32'Hfffffffe;
1434: data <= 32'H00000003;
1435: data <= 32'H00000006;
1436: data <= 32'H0000000a;
1437: data <= 32'H00000006;
1438: data <= 32'Hfffffffc;
1439: data <= 32'Hffffffff;
1440: data <= 32'Hfffffff8;
1441: data <= 32'Hfffffff9;
1442: data <= 32'Hfffffffd;
1443: data <= 32'Hfffffffe;
1444: data <= 32'Hfffffff7;
1445: data <= 32'Hfffffff6;
1446: data <= 32'Hfffffff0;
1447: data <= 32'Hffffffef;
1448: data <= 32'Hfffffff8;
1449: data <= 32'Hfffffff7;
1450: data <= 32'Hfffffff6;
1451: data <= 32'H00000001;
1452: data <= 32'H00000008;
1453: data <= 32'H00000007;
1454: data <= 32'H00000011;
1455: data <= 32'H0000000c;
1456: data <= 32'H00000000;
1457: data <= 32'Hfffffffe;
1458: data <= 32'Hfffffff8;
1459: data <= 32'Hffffffe8;
1460: data <= 32'Hffffffed;
1461: data <= 32'Hfffffff2;
1462: data <= 32'Hfffffffb;
1463: data <= 32'H00000007;
1464: data <= 32'H00000006;
1465: data <= 32'H00000007;
1466: data <= 32'H00000007;
1467: data <= 32'H00000004;
1468: data <= 32'H00000008;
1469: data <= 32'H0000000a;
1470: data <= 32'H0000000c;
1471: data <= 32'H0000000e;
1472: data <= 32'H00000009;
1473: data <= 32'H00000002;
1474: data <= 32'Hffffffff;
1475: data <= 32'Hfffffffc;
1476: data <= 32'Hfffffffa;
1477: data <= 32'H00000002;
1478: data <= 32'H00000002;
1479: data <= 32'H00000009;
1480: data <= 32'H0000000c;
1481: data <= 32'H0000000a;
1482: data <= 32'H00000004;
1483: data <= 32'H00000009;
1484: data <= 32'H00000006;
1485: data <= 32'H00000008;
1486: data <= 32'H00000005;
1487: data <= 32'H00000000;
1488: data <= 32'Hfffffffa;
1489: data <= 32'Hfffffffe;
1490: data <= 32'Hfffffffc;
1491: data <= 32'Hfffffffe;
1492: data <= 32'Hfffffffd;
1493: data <= 32'Hfffffffb;
1494: data <= 32'Hfffffff6;
1495: data <= 32'Hfffffff7;
1496: data <= 32'Hfffffff4;
1497: data <= 32'Hffffffef;
1498: data <= 32'Hffffffef;
1499: data <= 32'Hfffffff0;
1500: data <= 32'Hffffffee;
1501: data <= 32'Hffffffeb;
1502: data <= 32'Hffffffe8;
1503: data <= 32'Hffffffe8;
1504: data <= 32'Hffffffe7;
1505: data <= 32'Hffffffe5;
1506: data <= 32'Hffffffe8;
1507: data <= 32'Hffffffeb;
1508: data <= 32'Hffffffef;
1509: data <= 32'Hffffffee;
1510: data <= 32'Hfffffff4;
1511: data <= 32'Hfffffff7;
1512: data <= 32'Hfffffffd;
1513: data <= 32'Hfffffffd;
1514: data <= 32'H00000006;
1515: data <= 32'H00000009;
1516: data <= 32'H00000005;
1517: data <= 32'Hfffffffc;
1518: data <= 32'Hfffffff3;
1519: data <= 32'Hfffffff3;
1520: data <= 32'Hfffffff1;
1521: data <= 32'Hffffffed;
1522: data <= 32'Hfffffff7;
1523: data <= 32'Hffffffec;
1524: data <= 32'Hffffffe9;
1525: data <= 32'Hfffffff0;
1526: data <= 32'Hffffffef;
1527: data <= 32'Hffffffec;
1528: data <= 32'Hfffffff9;
1529: data <= 32'Hffffffff;
1530: data <= 32'Hfffffffd;
1531: data <= 32'H0000000c;
1532: data <= 32'H0000000e;
1533: data <= 32'H00000003;
1534: data <= 32'H00000004;
1535: data <= 32'H00000009;
1536: data <= 32'H0000000b;
1537: data <= 32'H00000003;
1538: data <= 32'H00000005;
1539: data <= 32'Hffffffff;
1540: data <= 32'H00000007;
1541: data <= 32'H00000002;
1542: data <= 32'H00000002;
1543: data <= 32'H00000006;
1544: data <= 32'H00000004;
1545: data <= 32'H00000005;
1546: data <= 32'H0000000a;
1547: data <= 32'H00000008;
1548: data <= 32'H00000004;
1549: data <= 32'H0000000a;
1550: data <= 32'H00000005;
1551: data <= 32'H0000000c;
1552: data <= 32'H00000009;
1553: data <= 32'H00000009;
1554: data <= 32'H00000005;
1555: data <= 32'H00000004;
1556: data <= 32'H00000001;
1557: data <= 32'Hffffffff;
1558: data <= 32'H00000001;
1559: data <= 32'Hffffffff;
1560: data <= 32'Hfffffffb;
1561: data <= 32'H00000003;
1562: data <= 32'H00000009;
1563: data <= 32'H00000003;
1564: data <= 32'H00000004;
1565: data <= 32'Hfffffffb;
1566: data <= 32'Hfffffff1;
1567: data <= 32'Hfffffff1;
1568: data <= 32'Hfffffff2;
1569: data <= 32'Hffffffef;
1570: data <= 32'Hffffffec;
1571: data <= 32'Hffffffed;
1572: data <= 32'Hffffffed;
1573: data <= 32'Hfffffff2;
1574: data <= 32'Hfffffff8;
1575: data <= 32'H00000001;
1576: data <= 32'H00000005;
1577: data <= 32'H00000002;
1578: data <= 32'H00000003;
1579: data <= 32'H00000006;
1580: data <= 32'H00000006;
1581: data <= 32'H00000009;
1582: data <= 32'H0000000b;
1583: data <= 32'H00000005;
1584: data <= 32'H00000000;
1585: data <= 32'Hfffffff9;
1586: data <= 32'Hfffffff8;
1587: data <= 32'Hfffffff3;
1588: data <= 32'Hfffffff7;
1589: data <= 32'H00000003;
1590: data <= 32'H00000009;
1591: data <= 32'H0000000c;
1592: data <= 32'H0000000c;
1593: data <= 32'H00000009;
1594: data <= 32'H00000005;
1595: data <= 32'H00000007;
1596: data <= 32'H0000000a;
1597: data <= 32'H00000011;
1598: data <= 32'H00000013;
1599: data <= 32'H0000000e;
1600: data <= 32'H00000008;
1601: data <= 32'Hffffffff;
1602: data <= 32'Hfffffffd;
1603: data <= 32'H00000000;
1604: data <= 32'H00000004;
1605: data <= 32'H00000009;
1606: data <= 32'H0000000e;
1607: data <= 32'H00000016;
1608: data <= 32'H00000013;
1609: data <= 32'H00000011;
1610: data <= 32'H0000000c;
1611: data <= 32'H0000000b;
1612: data <= 32'H00000008;
1613: data <= 32'H00000006;
1614: data <= 32'H00000000;
1615: data <= 32'Hfffffffb;
1616: data <= 32'Hfffffff9;
1617: data <= 32'Hfffffffe;
1618: data <= 32'Hfffffffe;
1619: data <= 32'Hffffffff;
1620: data <= 32'Hfffffffe;
1621: data <= 32'Hfffffffb;
1622: data <= 32'Hfffffffa;
1623: data <= 32'Hfffffff9;
1624: data <= 32'Hfffffff5;
1625: data <= 32'Hfffffff0;
1626: data <= 32'Hfffffff1;
1627: data <= 32'Hfffffff4;
1628: data <= 32'Hfffffff7;
1629: data <= 32'Hfffffff6;
1630: data <= 32'Hfffffff4;
1631: data <= 32'Hfffffff2;
1632: data <= 32'Hfffffff0;
1633: data <= 32'Hfffffff0;
1634: data <= 32'Hffffffea;
1635: data <= 32'Hffffffed;
1636: data <= 32'Hfffffff0;
1637: data <= 32'Hffffffed;
1638: data <= 32'Hfffffff5;
1639: data <= 32'Hfffffff4;
1640: data <= 32'Hfffffff6;
1641: data <= 32'H00000000;
1642: data <= 32'H00000009;
1643: data <= 32'H0000000f;
1644: data <= 32'H00000013;
1645: data <= 32'H0000000e;
1646: data <= 32'H00000009;
1647: data <= 32'H00000002;
1648: data <= 32'Hfffffffd;
1649: data <= 32'Hfffffffb;
1650: data <= 32'Hfffffff9;
1651: data <= 32'Hfffffff7;
1652: data <= 32'Hfffffff4;
1653: data <= 32'Hfffffff4;
1654: data <= 32'Hfffffff0;
1655: data <= 32'Hfffffff0;
1656: data <= 32'Hfffffff3;
1657: data <= 32'Hfffffff7;
1658: data <= 32'Hfffffff3;
1659: data <= 32'Hffffffff;
1660: data <= 32'H0000000a;
1661: data <= 32'H00000006;
1662: data <= 32'H00000008;
1663: data <= 32'H0000000e;
1664: data <= 32'H0000000e;
1665: data <= 32'H0000000d;
1666: data <= 32'H00000013;
1667: data <= 32'H00000014;
1668: data <= 32'H00000012;
1669: data <= 32'H00000010;
1670: data <= 32'H0000000f;
1671: data <= 32'H00000013;
1672: data <= 32'H0000000f;
1673: data <= 32'H00000011;
1674: data <= 32'H0000000f;
1675: data <= 32'H00000016;
1676: data <= 32'H0000000f;
1677: data <= 32'H00000012;
1678: data <= 32'H00000016;
1679: data <= 32'H00000017;
1680: data <= 32'H00000015;
1681: data <= 32'H00000017;
1682: data <= 32'H0000000f;
1683: data <= 32'H0000000e;
1684: data <= 32'H00000011;
1685: data <= 32'H0000000c;
1686: data <= 32'H0000000f;
1687: data <= 32'H00000010;
1688: data <= 32'H0000000e;
1689: data <= 32'H0000000f;
1690: data <= 32'H00000016;
1691: data <= 32'H0000000f;
1692: data <= 32'H00000008;
1693: data <= 32'H00000003;
1694: data <= 32'Hfffffffe;
1695: data <= 32'Hfffffffb;
1696: data <= 32'Hfffffffc;
1697: data <= 32'Hfffffff8;
1698: data <= 32'Hfffffffc;
1699: data <= 32'H00000004;
1700: data <= 32'H0000000d;
1701: data <= 32'H00000016;
1702: data <= 32'H0000001c;
1703: data <= 32'H0000001a;
1704: data <= 32'H00000019;
1705: data <= 32'H00000014;
1706: data <= 32'H0000000e;
1707: data <= 32'H0000000f;
1708: data <= 32'H0000000c;
1709: data <= 32'H00000008;
1710: data <= 32'H0000000b;
1711: data <= 32'H00000005;
1712: data <= 32'H00000002;
1713: data <= 32'Hfffffffe;
1714: data <= 32'Hfffffff7;
1715: data <= 32'Hfffffff7;
1716: data <= 32'Hfffffffc;
1717: data <= 32'H00000004;
1718: data <= 32'H00000007;
1719: data <= 32'H0000000b;
1720: data <= 32'H00000006;
1721: data <= 32'H00000005;
1722: data <= 32'H00000001;
1723: data <= 32'H0000000a;
1724: data <= 32'H0000000c;
1725: data <= 32'H00000010;
1726: data <= 32'H0000000d;
1727: data <= 32'H00000009;
1728: data <= 32'H00000005;
1729: data <= 32'Hfffffffe;
1730: data <= 32'H00000002;
1731: data <= 32'H0000000a;
1732: data <= 32'H0000000a;
1733: data <= 32'H0000000b;
1734: data <= 32'H00000011;
1735: data <= 32'H00000014;
1736: data <= 32'H00000013;
1737: data <= 32'H0000000f;
1738: data <= 32'H0000000f;
1739: data <= 32'H0000000a;
1740: data <= 32'H00000005;
1741: data <= 32'Hffffffff;
1742: data <= 32'Hfffffff8;
1743: data <= 32'Hfffffff6;
1744: data <= 32'Hfffffff6;
1745: data <= 32'Hfffffff9;
1746: data <= 32'Hfffffffb;
1747: data <= 32'Hfffffffa;
1748: data <= 32'Hfffffff9;
1749: data <= 32'Hfffffff8;
1750: data <= 32'Hfffffff7;
1751: data <= 32'Hffffffef;
1752: data <= 32'Hffffffee;
1753: data <= 32'Hffffffea;
1754: data <= 32'Hffffffee;
1755: data <= 32'Hfffffff2;
1756: data <= 32'Hfffffffa;
1757: data <= 32'Hfffffffc;
1758: data <= 32'Hfffffffd;
1759: data <= 32'H00000001;
1760: data <= 32'Hffffffff;
1761: data <= 32'Hffffffff;
1762: data <= 32'Hfffffff7;
1763: data <= 32'Hfffffff3;
1764: data <= 32'Hfffffff6;
1765: data <= 32'Hfffffff4;
1766: data <= 32'Hfffffff9;
1767: data <= 32'Hfffffffa;
1768: data <= 32'Hfffffffa;
1769: data <= 32'Hfffffffd;
1770: data <= 32'H00000005;
1771: data <= 32'H00000009;
1772: data <= 32'H00000013;
1773: data <= 32'H00000014;
1774: data <= 32'H0000000f;
1775: data <= 32'H00000010;
1776: data <= 32'H0000000d;
1777: data <= 32'H0000000c;
1778: data <= 32'H00000009;
1779: data <= 32'H00000004;
1780: data <= 32'H00000002;
1781: data <= 32'H00000001;
1782: data <= 32'Hfffffffb;
1783: data <= 32'Hfffffffa;
1784: data <= 32'Hfffffffb;
1785: data <= 32'Hfffffffa;
1786: data <= 32'Hfffffffc;
1787: data <= 32'Hfffffffb;
1788: data <= 32'Hfffffffd;
1789: data <= 32'H00000001;
1790: data <= 32'H00000008;
1791: data <= 32'H00000008;
1792: data <= 32'H0000000c;
1793: data <= 32'Hfffffffd;
1794: data <= 32'H00000000;
1795: data <= 32'H00000002;
1796: data <= 32'H00000002;
1797: data <= 32'H00000002;
1798: data <= 32'Hfffffffd;
1799: data <= 32'H00000002;
1800: data <= 32'H00000001;
1801: data <= 32'H00000007;
1802: data <= 32'H00000002;
1803: data <= 32'H00000005;
1804: data <= 32'H00000006;
1805: data <= 32'H00000009;
1806: data <= 32'H00000005;
1807: data <= 32'H0000000c;
1808: data <= 32'H00000006;
1809: data <= 32'H00000003;
1810: data <= 32'H00000005;
1811: data <= 32'H00000004;
1812: data <= 32'H00000007;
1813: data <= 32'H0000000a;
1814: data <= 32'H00000007;
1815: data <= 32'H00000004;
1816: data <= 32'H0000000a;
1817: data <= 32'H00000003;
1818: data <= 32'H00000007;
1819: data <= 32'H00000003;
1820: data <= 32'H00000000;
1821: data <= 32'Hfffffff5;
1822: data <= 32'Hfffffffa;
1823: data <= 32'Hfffffff4;
1824: data <= 32'Hfffffff9;
1825: data <= 32'H00000002;
1826: data <= 32'H00000007;
1827: data <= 32'H0000000c;
1828: data <= 32'H00000014;
1829: data <= 32'H00000012;
1830: data <= 32'H00000012;
1831: data <= 32'H0000000f;
1832: data <= 32'H0000000c;
1833: data <= 32'H00000008;
1834: data <= 32'H00000004;
1835: data <= 32'Hfffffff9;
1836: data <= 32'Hfffffff8;
1837: data <= 32'Hfffffff7;
1838: data <= 32'Hfffffff3;
1839: data <= 32'Hfffffff0;
1840: data <= 32'Hffffffe9;
1841: data <= 32'Hffffffe3;
1842: data <= 32'Hffffffe1;
1843: data <= 32'Hffffffeb;
1844: data <= 32'Hffffffeb;
1845: data <= 32'Hfffffff5;
1846: data <= 32'Hfffffff2;
1847: data <= 32'Hfffffff2;
1848: data <= 32'Hffffffea;
1849: data <= 32'Hffffffeb;
1850: data <= 32'Hffffffec;
1851: data <= 32'Hfffffff1;
1852: data <= 32'Hfffffff2;
1853: data <= 32'Hfffffffb;
1854: data <= 32'Hfffffffc;
1855: data <= 32'Hfffffffb;
1856: data <= 32'Hfffffffc;
1857: data <= 32'Hfffffffd;
1858: data <= 32'H00000004;
1859: data <= 32'H0000000a;
1860: data <= 32'H0000000c;
1861: data <= 32'H0000000e;
1862: data <= 32'H00000011;
1863: data <= 32'H00000010;
1864: data <= 32'H0000000c;
1865: data <= 32'H00000008;
1866: data <= 32'H00000004;
1867: data <= 32'H00000000;
1868: data <= 32'Hfffffff7;
1869: data <= 32'Hfffffff0;
1870: data <= 32'Hffffffe6;
1871: data <= 32'Hffffffe6;
1872: data <= 32'Hffffffeb;
1873: data <= 32'Hffffffe8;
1874: data <= 32'Hffffffeb;
1875: data <= 32'Hffffffeb;
1876: data <= 32'Hffffffec;
1877: data <= 32'Hffffffec;
1878: data <= 32'Hffffffee;
1879: data <= 32'Hffffffe3;
1880: data <= 32'Hffffffe3;
1881: data <= 32'Hffffffe3;
1882: data <= 32'Hffffffe4;
1883: data <= 32'Hffffffe8;
1884: data <= 32'Hfffffff0;
1885: data <= 32'Hfffffff6;
1886: data <= 32'Hfffffffc;
1887: data <= 32'H00000000;
1888: data <= 32'H00000001;
1889: data <= 32'H00000002;
1890: data <= 32'H00000001;
1891: data <= 32'Hfffffffb;
1892: data <= 32'Hfffffff8;
1893: data <= 32'Hfffffff8;
1894: data <= 32'Hfffffff9;
1895: data <= 32'Hfffffff6;
1896: data <= 32'Hfffffffa;
1897: data <= 32'Hfffffff3;
1898: data <= 32'Hfffffff1;
1899: data <= 32'Hfffffff5;
1900: data <= 32'Hfffffff9;
1901: data <= 32'Hfffffffa;
1902: data <= 32'Hfffffffc;
1903: data <= 32'Hfffffffa;
1904: data <= 32'Hfffffffb;
1905: data <= 32'H00000001;
1906: data <= 32'Hfffffffe;
1907: data <= 32'H00000000;
1908: data <= 32'H00000000;
1909: data <= 32'Hfffffffc;
1910: data <= 32'Hfffffffa;
1911: data <= 32'Hfffffff1;
1912: data <= 32'Hffffffef;
1913: data <= 32'Hffffffef;
1914: data <= 32'Hfffffff3;
1915: data <= 32'Hffffffea;
1916: data <= 32'Hfffffff0;
1917: data <= 32'Hffffffee;
1918: data <= 32'Hffffffed;
1919: data <= 32'Hffffffec;
1920: data <= 32'Hfffffff4;
1921: data <= 32'H00000000;
1922: data <= 32'Hfffffffe;
1923: data <= 32'H00000003;
1924: data <= 32'Hfffffffe;
1925: data <= 32'H00000005;
1926: data <= 32'Hffffffff;
1927: data <= 32'H00000000;
1928: data <= 32'H00000006;
1929: data <= 32'H00000009;
1930: data <= 32'H00000004;
1931: data <= 32'H0000000b;
1932: data <= 32'H0000000b;
1933: data <= 32'H00000009;
1934: data <= 32'H0000000e;
1935: data <= 32'H0000000b;
1936: data <= 32'H00000007;
1937: data <= 32'H00000003;
1938: data <= 32'H00000006;
1939: data <= 32'H0000000b;
1940: data <= 32'H0000000d;
1941: data <= 32'H00000011;
1942: data <= 32'H0000000b;
1943: data <= 32'H00000006;
1944: data <= 32'H0000000d;
1945: data <= 32'H0000000a;
1946: data <= 32'H0000000a;
1947: data <= 32'H00000005;
1948: data <= 32'Hfffffffd;
1949: data <= 32'Hfffffffb;
1950: data <= 32'H00000003;
1951: data <= 32'H00000006;
1952: data <= 32'H00000011;
1953: data <= 32'H00000013;
1954: data <= 32'H00000015;
1955: data <= 32'H00000014;
1956: data <= 32'H00000013;
1957: data <= 32'H00000010;
1958: data <= 32'H0000000f;
1959: data <= 32'H00000003;
1960: data <= 32'H00000000;
1961: data <= 32'Hfffffffd;
1962: data <= 32'Hfffffff3;
1963: data <= 32'Hfffffff1;
1964: data <= 32'Hffffffe9;
1965: data <= 32'Hffffffe7;
1966: data <= 32'Hffffffe3;
1967: data <= 32'Hffffffe0;
1968: data <= 32'Hffffffdf;
1969: data <= 32'Hffffffe1;
1970: data <= 32'Hffffffe0;
1971: data <= 32'Hffffffee;
1972: data <= 32'Hfffffff0;
1973: data <= 32'Hfffffff2;
1974: data <= 32'Hffffffed;
1975: data <= 32'Hffffffe8;
1976: data <= 32'Hffffffdf;
1977: data <= 32'Hffffffe4;
1978: data <= 32'Hffffffe4;
1979: data <= 32'Hffffffea;
1980: data <= 32'Hfffffff0;
1981: data <= 32'Hfffffffc;
1982: data <= 32'H00000005;
1983: data <= 32'H00000006;
1984: data <= 32'H0000000b;
1985: data <= 32'H00000015;
1986: data <= 32'H00000015;
1987: data <= 32'H00000018;
1988: data <= 32'H0000001b;
1989: data <= 32'H00000019;
1990: data <= 32'H0000001b;
1991: data <= 32'H0000001a;
1992: data <= 32'H00000014;
1993: data <= 32'H0000000e;
1994: data <= 32'H00000009;
1995: data <= 32'H00000007;
1996: data <= 32'Hfffffffe;
1997: data <= 32'Hfffffff2;
1998: data <= 32'Hffffffef;
1999: data <= 32'Hffffffef;
2000: data <= 32'Hfffffff3;
2001: data <= 32'Hfffffff3;
2002: data <= 32'Hfffffffb;
2003: data <= 32'Hfffffffa;
2004: data <= 32'Hfffffff9;
2005: data <= 32'Hfffffff8;
2006: data <= 32'Hfffffff8;
2007: data <= 32'Hfffffff0;
2008: data <= 32'Hffffffef;
2009: data <= 32'Hfffffff2;
2010: data <= 32'Hfffffff0;
2011: data <= 32'Hfffffff3;
2012: data <= 32'Hfffffffe;
2013: data <= 32'H00000005;
2014: data <= 32'H00000008;
2015: data <= 32'H0000000a;
2016: data <= 32'H00000008;
2017: data <= 32'H0000000d;
2018: data <= 32'H0000000e;
2019: data <= 32'H00000007;
2020: data <= 32'H00000007;
2021: data <= 32'H00000004;
2022: data <= 32'Hfffffffe;
2023: data <= 32'Hfffffffb;
2024: data <= 32'Hfffffff8;
2025: data <= 32'Hffffffef;
2026: data <= 32'Hffffffec;
2027: data <= 32'Hffffffeb;
2028: data <= 32'Hfffffff2;
2029: data <= 32'Hffffffef;
2030: data <= 32'Hffffffee;
2031: data <= 32'Hffffffeb;
2032: data <= 32'Hffffffe7;
2033: data <= 32'Hffffffe7;
2034: data <= 32'Hfffffff1;
2035: data <= 32'Hfffffff5;
2036: data <= 32'Hfffffffb;
2037: data <= 32'H00000003;
2038: data <= 32'H00000002;
2039: data <= 32'Hfffffff7;
2040: data <= 32'Hfffffff0;
2041: data <= 32'Hffffffeb;
2042: data <= 32'Hffffffee;
2043: data <= 32'Hfffffff0;
2044: data <= 32'Hfffffff6;
2045: data <= 32'Hfffffff2;
2046: data <= 32'Hffffffee;
2047: data <= 32'Hffffffe5;
2048: data <= 32'Hffffffee;
2049: data <= 32'H00000006;
2050: data <= 32'Hfffffffd;
2051: data <= 32'Hffffffff;
2052: data <= 32'H00000000;
2053: data <= 32'H00000001;
2054: data <= 32'H00000003;
2055: data <= 32'H00000004;
2056: data <= 32'H00000009;
2057: data <= 32'H00000007;
2058: data <= 32'H0000000a;
2059: data <= 32'H0000000c;
2060: data <= 32'H0000000d;
2061: data <= 32'H0000000d;
2062: data <= 32'H0000000f;
2063: data <= 32'H0000000a;
2064: data <= 32'H00000007;
2065: data <= 32'H00000007;
2066: data <= 32'H00000007;
2067: data <= 32'H0000000a;
2068: data <= 32'H00000008;
2069: data <= 32'H00000008;
2070: data <= 32'H00000000;
2071: data <= 32'Hfffffffe;
2072: data <= 32'H00000002;
2073: data <= 32'Hffffffff;
2074: data <= 32'Hfffffffb;
2075: data <= 32'Hfffffff4;
2076: data <= 32'Hfffffff7;
2077: data <= 32'Hfffffffe;
2078: data <= 32'H0000000a;
2079: data <= 32'H00000012;
2080: data <= 32'H00000011;
2081: data <= 32'H0000000d;
2082: data <= 32'H0000000f;
2083: data <= 32'H0000000e;
2084: data <= 32'H0000000d;
2085: data <= 32'H0000000b;
2086: data <= 32'H00000003;
2087: data <= 32'Hffffffff;
2088: data <= 32'Hfffffffa;
2089: data <= 32'Hfffffffa;
2090: data <= 32'Hfffffff7;
2091: data <= 32'Hffffffef;
2092: data <= 32'Hffffffe5;
2093: data <= 32'Hffffffe3;
2094: data <= 32'Hffffffe9;
2095: data <= 32'Hffffffeb;
2096: data <= 32'Hffffffec;
2097: data <= 32'Hfffffff3;
2098: data <= 32'Hfffffff6;
2099: data <= 32'Hfffffffa;
2100: data <= 32'Hfffffffd;
2101: data <= 32'Hfffffffc;
2102: data <= 32'Hffffffec;
2103: data <= 32'Hffffffea;
2104: data <= 32'Hffffffe4;
2105: data <= 32'Hffffffe0;
2106: data <= 32'Hffffffe6;
2107: data <= 32'Hffffffec;
2108: data <= 32'Hfffffff7;
2109: data <= 32'H00000003;
2110: data <= 32'H0000000b;
2111: data <= 32'H00000011;
2112: data <= 32'H00000015;
2113: data <= 32'H00000017;
2114: data <= 32'H0000001c;
2115: data <= 32'H0000001a;
2116: data <= 32'H00000017;
2117: data <= 32'H00000019;
2118: data <= 32'H00000017;
2119: data <= 32'H00000013;
2120: data <= 32'H00000011;
2121: data <= 32'H00000008;
2122: data <= 32'H00000002;
2123: data <= 32'H00000004;
2124: data <= 32'Hfffffffe;
2125: data <= 32'Hfffffff3;
2126: data <= 32'Hfffffff5;
2127: data <= 32'Hfffffff0;
2128: data <= 32'Hfffffff6;
2129: data <= 32'Hfffffff9;
2130: data <= 32'Hfffffffb;
2131: data <= 32'Hfffffffa;
2132: data <= 32'Hfffffffa;
2133: data <= 32'Hfffffff4;
2134: data <= 32'Hfffffff0;
2135: data <= 32'Hffffffee;
2136: data <= 32'Hffffffea;
2137: data <= 32'Hffffffea;
2138: data <= 32'Hffffffec;
2139: data <= 32'Hfffffff1;
2140: data <= 32'Hfffffff8;
2141: data <= 32'H00000000;
2142: data <= 32'H00000002;
2143: data <= 32'H00000000;
2144: data <= 32'H00000008;
2145: data <= 32'H00000007;
2146: data <= 32'H00000004;
2147: data <= 32'Hfffffffd;
2148: data <= 32'Hfffffffa;
2149: data <= 32'Hffffffff;
2150: data <= 32'Hfffffffa;
2151: data <= 32'Hfffffff9;
2152: data <= 32'Hfffffff2;
2153: data <= 32'Hffffffeb;
2154: data <= 32'Hffffffe9;
2155: data <= 32'Hffffffe8;
2156: data <= 32'Hffffffec;
2157: data <= 32'Hfffffff0;
2158: data <= 32'Hfffffff0;
2159: data <= 32'Hffffffe8;
2160: data <= 32'Hffffffe7;
2161: data <= 32'Hffffffdf;
2162: data <= 32'Hffffffe4;
2163: data <= 32'Hffffffe7;
2164: data <= 32'Hffffffec;
2165: data <= 32'Hfffffff1;
2166: data <= 32'Hfffffff8;
2167: data <= 32'Hfffffff5;
2168: data <= 32'Hfffffff4;
2169: data <= 32'Hfffffff1;
2170: data <= 32'Hffffffea;
2171: data <= 32'Hffffffe9;
2172: data <= 32'Hfffffff3;
2173: data <= 32'Hfffffff0;
2174: data <= 32'Hffffffee;
2175: data <= 32'Hffffffec;
2176: data <= 32'Hffffffec;
2177: data <= 32'Hfffffffd;
2178: data <= 32'Hfffffff8;
2179: data <= 32'Hfffffff6;
2180: data <= 32'Hfffffffe;
2181: data <= 32'Hfffffffa;
2182: data <= 32'Hfffffffd;
2183: data <= 32'Hfffffffe;
2184: data <= 32'H00000000;
2185: data <= 32'Hfffffffc;
2186: data <= 32'H00000003;
2187: data <= 32'H00000002;
2188: data <= 32'H00000003;
2189: data <= 32'H00000003;
2190: data <= 32'H00000006;
2191: data <= 32'H00000000;
2192: data <= 32'H00000000;
2193: data <= 32'H00000001;
2194: data <= 32'Hfffffffd;
2195: data <= 32'Hffffffff;
2196: data <= 32'Hfffffff7;
2197: data <= 32'Hfffffff4;
2198: data <= 32'Hffffffed;
2199: data <= 32'Hffffffee;
2200: data <= 32'Hffffffec;
2201: data <= 32'Hfffffff2;
2202: data <= 32'Hfffffff3;
2203: data <= 32'Hfffffff3;
2204: data <= 32'Hfffffff6;
2205: data <= 32'H00000006;
2206: data <= 32'H00000006;
2207: data <= 32'H0000000e;
2208: data <= 32'H0000000b;
2209: data <= 32'H00000009;
2210: data <= 32'H0000000a;
2211: data <= 32'H0000000c;
2212: data <= 32'H0000000d;
2213: data <= 32'H00000008;
2214: data <= 32'H00000000;
2215: data <= 32'H00000002;
2216: data <= 32'H00000000;
2217: data <= 32'Hfffffffb;
2218: data <= 32'Hfffffff6;
2219: data <= 32'Hfffffff0;
2220: data <= 32'Hffffffe8;
2221: data <= 32'Hffffffe9;
2222: data <= 32'Hfffffff2;
2223: data <= 32'Hfffffff5;
2224: data <= 32'Hfffffffb;
2225: data <= 32'Hfffffffa;
2226: data <= 32'H00000000;
2227: data <= 32'H00000001;
2228: data <= 32'H00000001;
2229: data <= 32'Hfffffff3;
2230: data <= 32'Hffffffeb;
2231: data <= 32'Hffffffe3;
2232: data <= 32'Hffffffe3;
2233: data <= 32'Hffffffe0;
2234: data <= 32'Hffffffe3;
2235: data <= 32'Hffffffea;
2236: data <= 32'Hfffffff8;
2237: data <= 32'H00000000;
2238: data <= 32'H0000000a;
2239: data <= 32'H0000000c;
2240: data <= 32'H0000000a;
2241: data <= 32'H00000010;
2242: data <= 32'H0000000f;
2243: data <= 32'H0000000f;
2244: data <= 32'H0000000c;
2245: data <= 32'H0000000a;
2246: data <= 32'H0000000b;
2247: data <= 32'H00000007;
2248: data <= 32'H00000004;
2249: data <= 32'H00000002;
2250: data <= 32'H00000002;
2251: data <= 32'H00000000;
2252: data <= 32'H00000000;
2253: data <= 32'Hfffffffc;
2254: data <= 32'Hfffffff6;
2255: data <= 32'Hfffffff6;
2256: data <= 32'Hfffffff5;
2257: data <= 32'Hfffffff4;
2258: data <= 32'Hfffffff2;
2259: data <= 32'Hfffffff2;
2260: data <= 32'Hffffffea;
2261: data <= 32'Hffffffeb;
2262: data <= 32'Hffffffe7;
2263: data <= 32'Hffffffe4;
2264: data <= 32'Hffffffe3;
2265: data <= 32'Hffffffe1;
2266: data <= 32'Hffffffe7;
2267: data <= 32'Hffffffec;
2268: data <= 32'Hfffffff2;
2269: data <= 32'Hfffffff3;
2270: data <= 32'Hfffffff6;
2271: data <= 32'Hfffffff9;
2272: data <= 32'Hffffffff;
2273: data <= 32'Hffffffff;
2274: data <= 32'Hfffffff9;
2275: data <= 32'Hfffffffc;
2276: data <= 32'Hfffffff8;
2277: data <= 32'Hfffffff9;
2278: data <= 32'Hfffffffc;
2279: data <= 32'H00000002;
2280: data <= 32'Hfffffffe;
2281: data <= 32'H00000004;
2282: data <= 32'H00000003;
2283: data <= 32'H00000000;
2284: data <= 32'H00000001;
2285: data <= 32'H00000000;
2286: data <= 32'Hfffffffe;
2287: data <= 32'Hfffffffc;
2288: data <= 32'Hfffffff6;
2289: data <= 32'Hffffffed;
2290: data <= 32'Hffffffec;
2291: data <= 32'Hffffffe8;
2292: data <= 32'Hffffffe2;
2293: data <= 32'Hffffffdf;
2294: data <= 32'Hffffffdb;
2295: data <= 32'Hffffffdd;
2296: data <= 32'Hffffffe0;
2297: data <= 32'Hffffffe4;
2298: data <= 32'Hffffffe0;
2299: data <= 32'Hffffffe0;
2300: data <= 32'Hffffffdd;
2301: data <= 32'Hffffffdd;
2302: data <= 32'Hffffffe2;
2303: data <= 32'Hffffffe3;
2304: data <= 32'Hffffffe1;
2305: data <= 32'Hffffffff;
2306: data <= 32'H00000001;
2307: data <= 32'H00000000;
2308: data <= 32'H00000005;
2309: data <= 32'Hfffffffe;
2310: data <= 32'H00000002;
2311: data <= 32'H00000003;
2312: data <= 32'H00000000;
2313: data <= 32'H00000000;
2314: data <= 32'H00000001;
2315: data <= 32'H00000003;
2316: data <= 32'H00000000;
2317: data <= 32'H00000001;
2318: data <= 32'Hffffffff;
2319: data <= 32'H00000001;
2320: data <= 32'Hfffffffe;
2321: data <= 32'Hfffffffd;
2322: data <= 32'Hfffffff9;
2323: data <= 32'Hfffffffc;
2324: data <= 32'Hfffffffb;
2325: data <= 32'Hfffffff0;
2326: data <= 32'Hffffffea;
2327: data <= 32'Hffffffec;
2328: data <= 32'Hffffffea;
2329: data <= 32'Hfffffff1;
2330: data <= 32'Hfffffff5;
2331: data <= 32'Hfffffff4;
2332: data <= 32'Hfffffffc;
2333: data <= 32'H00000000;
2334: data <= 32'H00000001;
2335: data <= 32'H00000007;
2336: data <= 32'H00000005;
2337: data <= 32'H00000005;
2338: data <= 32'H00000008;
2339: data <= 32'H00000008;
2340: data <= 32'H00000009;
2341: data <= 32'H00000003;
2342: data <= 32'Hfffffffe;
2343: data <= 32'Hffffffff;
2344: data <= 32'Hfffffffd;
2345: data <= 32'Hfffffff9;
2346: data <= 32'Hfffffff4;
2347: data <= 32'Hfffffff0;
2348: data <= 32'Hfffffff2;
2349: data <= 32'Hfffffff3;
2350: data <= 32'Hfffffffc;
2351: data <= 32'Hfffffffe;
2352: data <= 32'H00000003;
2353: data <= 32'H00000002;
2354: data <= 32'H00000003;
2355: data <= 32'H00000001;
2356: data <= 32'Hfffffffb;
2357: data <= 32'Hfffffff0;
2358: data <= 32'Hffffffeb;
2359: data <= 32'Hffffffeb;
2360: data <= 32'Hffffffe7;
2361: data <= 32'Hffffffe3;
2362: data <= 32'Hffffffe8;
2363: data <= 32'Hffffffe9;
2364: data <= 32'Hfffffff5;
2365: data <= 32'Hffffffff;
2366: data <= 32'H00000001;
2367: data <= 32'H00000001;
2368: data <= 32'H00000006;
2369: data <= 32'H00000002;
2370: data <= 32'H00000004;
2371: data <= 32'H00000006;
2372: data <= 32'H00000000;
2373: data <= 32'Hffffffff;
2374: data <= 32'H00000005;
2375: data <= 32'H00000002;
2376: data <= 32'H00000003;
2377: data <= 32'H00000003;
2378: data <= 32'H00000000;
2379: data <= 32'Hffffffff;
2380: data <= 32'H00000001;
2381: data <= 32'Hfffffffa;
2382: data <= 32'Hfffffff7;
2383: data <= 32'Hfffffff9;
2384: data <= 32'Hfffffff7;
2385: data <= 32'Hfffffff7;
2386: data <= 32'Hfffffff1;
2387: data <= 32'Hfffffff2;
2388: data <= 32'Hffffffee;
2389: data <= 32'Hffffffeb;
2390: data <= 32'Hffffffe9;
2391: data <= 32'Hffffffe6;
2392: data <= 32'Hffffffe6;
2393: data <= 32'Hffffffe6;
2394: data <= 32'Hffffffed;
2395: data <= 32'Hfffffff1;
2396: data <= 32'Hfffffff4;
2397: data <= 32'Hfffffff5;
2398: data <= 32'Hfffffff8;
2399: data <= 32'Hfffffff8;
2400: data <= 32'Hfffffffc;
2401: data <= 32'Hfffffffd;
2402: data <= 32'Hfffffff7;
2403: data <= 32'H00000001;
2404: data <= 32'Hffffffff;
2405: data <= 32'Hfffffffb;
2406: data <= 32'H00000004;
2407: data <= 32'H0000000a;
2408: data <= 32'H0000000e;
2409: data <= 32'H00000019;
2410: data <= 32'H0000001b;
2411: data <= 32'H0000001a;
2412: data <= 32'H0000001a;
2413: data <= 32'H0000001d;
2414: data <= 32'H0000000d;
2415: data <= 32'H00000008;
2416: data <= 32'Hfffffffc;
2417: data <= 32'Hfffffff5;
2418: data <= 32'Hfffffff7;
2419: data <= 32'Hfffffff3;
2420: data <= 32'Hffffffed;
2421: data <= 32'Hffffffe2;
2422: data <= 32'Hffffffd4;
2423: data <= 32'Hffffffd1;
2424: data <= 32'Hffffffd9;
2425: data <= 32'Hffffffdd;
2426: data <= 32'Hffffffe3;
2427: data <= 32'Hffffffea;
2428: data <= 32'Hffffffe7;
2429: data <= 32'Hffffffea;
2430: data <= 32'Hffffffe9;
2431: data <= 32'Hffffffeb;
2432: data <= 32'Hffffffe7;
2433: data <= 32'Hfffffff0;
2434: data <= 32'Hfffffff6;
2435: data <= 32'Hfffffff6;
2436: data <= 32'Hfffffff4;
2437: data <= 32'Hfffffff5;
2438: data <= 32'Hfffffff6;
2439: data <= 32'Hfffffff7;
2440: data <= 32'Hfffffff2;
2441: data <= 32'Hfffffff8;
2442: data <= 32'Hfffffff1;
2443: data <= 32'Hfffffff2;
2444: data <= 32'Hffffffee;
2445: data <= 32'Hffffffef;
2446: data <= 32'Hffffffeb;
2447: data <= 32'Hfffffff3;
2448: data <= 32'Hffffffed;
2449: data <= 32'Hffffffef;
2450: data <= 32'Hfffffff0;
2451: data <= 32'Hfffffff0;
2452: data <= 32'Hfffffff5;
2453: data <= 32'Hffffffe5;
2454: data <= 32'Hffffffdc;
2455: data <= 32'Hffffffdc;
2456: data <= 32'Hffffffe3;
2457: data <= 32'Hffffffe8;
2458: data <= 32'Hffffffee;
2459: data <= 32'Hffffffee;
2460: data <= 32'Hfffffff1;
2461: data <= 32'Hfffffff4;
2462: data <= 32'Hfffffffa;
2463: data <= 32'Hfffffff5;
2464: data <= 32'Hfffffff7;
2465: data <= 32'Hfffffff7;
2466: data <= 32'Hfffffffd;
2467: data <= 32'Hfffffffa;
2468: data <= 32'Hfffffffc;
2469: data <= 32'Hfffffff2;
2470: data <= 32'Hffffffed;
2471: data <= 32'Hffffffeb;
2472: data <= 32'Hffffffea;
2473: data <= 32'Hffffffe6;
2474: data <= 32'Hffffffe6;
2475: data <= 32'Hffffffe2;
2476: data <= 32'Hffffffe6;
2477: data <= 32'Hffffffed;
2478: data <= 32'Hffffffed;
2479: data <= 32'Hfffffff5;
2480: data <= 32'Hfffffffb;
2481: data <= 32'Hfffffff3;
2482: data <= 32'Hffffffeb;
2483: data <= 32'Hffffffea;
2484: data <= 32'Hffffffe3;
2485: data <= 32'Hffffffe5;
2486: data <= 32'Hffffffe4;
2487: data <= 32'Hffffffe3;
2488: data <= 32'Hffffffde;
2489: data <= 32'Hffffffdb;
2490: data <= 32'Hffffffde;
2491: data <= 32'Hffffffe3;
2492: data <= 32'Hffffffe8;
2493: data <= 32'Hffffffe8;
2494: data <= 32'Hffffffee;
2495: data <= 32'Hffffffed;
2496: data <= 32'Hffffffec;
2497: data <= 32'Hffffffef;
2498: data <= 32'Hffffffed;
2499: data <= 32'Hffffffed;
2500: data <= 32'Hfffffff3;
2501: data <= 32'Hffffffef;
2502: data <= 32'Hfffffff8;
2503: data <= 32'Hfffffff5;
2504: data <= 32'Hfffffff0;
2505: data <= 32'Hffffffeb;
2506: data <= 32'Hffffffee;
2507: data <= 32'Hffffffea;
2508: data <= 32'Hffffffee;
2509: data <= 32'Hffffffec;
2510: data <= 32'Hffffffe8;
2511: data <= 32'Hffffffea;
2512: data <= 32'Hffffffea;
2513: data <= 32'Hffffffe7;
2514: data <= 32'Hffffffe8;
2515: data <= 32'Hffffffe7;
2516: data <= 32'Hffffffe2;
2517: data <= 32'Hffffffe1;
2518: data <= 32'Hffffffe4;
2519: data <= 32'Hffffffdb;
2520: data <= 32'Hffffffe1;
2521: data <= 32'Hffffffe2;
2522: data <= 32'Hffffffe9;
2523: data <= 32'Hffffffea;
2524: data <= 32'Hffffffef;
2525: data <= 32'Hffffffef;
2526: data <= 32'Hfffffff1;
2527: data <= 32'Hfffffff2;
2528: data <= 32'Hffffffee;
2529: data <= 32'Hfffffff1;
2530: data <= 32'Hffffffeb;
2531: data <= 32'Hffffffee;
2532: data <= 32'Hffffffef;
2533: data <= 32'Hfffffff4;
2534: data <= 32'Hfffffff8;
2535: data <= 32'Hfffffffe;
2536: data <= 32'H00000006;
2537: data <= 32'H0000000c;
2538: data <= 32'H00000008;
2539: data <= 32'H0000000c;
2540: data <= 32'H0000000a;
2541: data <= 32'H00000013;
2542: data <= 32'H00000012;
2543: data <= 32'H0000000b;
2544: data <= 32'Hfffffff9;
2545: data <= 32'Hffffffed;
2546: data <= 32'Hffffffe5;
2547: data <= 32'Hffffffe3;
2548: data <= 32'Hffffffeb;
2549: data <= 32'Hffffffe4;
2550: data <= 32'Hffffffdb;
2551: data <= 32'Hffffffcf;
2552: data <= 32'Hffffffcc;
2553: data <= 32'Hffffffd3;
2554: data <= 32'Hffffffe1;
2555: data <= 32'Hffffffeb;
2556: data <= 32'Hfffffff7;
2557: data <= 32'Hfffffffb;
2558: data <= 32'Hfffffffc;
2559: data <= 32'Hfffffff7;
2560: data <= 32'Hffffffed;
2561: data <= 32'Hfffffff6;
2562: data <= 32'Hfffffff9;
2563: data <= 32'Hfffffff9;
2564: data <= 32'Hfffffff5;
2565: data <= 32'Hfffffffb;
2566: data <= 32'Hfffffffb;
2567: data <= 32'Hfffffff9;
2568: data <= 32'Hfffffffd;
2569: data <= 32'H00000001;
2570: data <= 32'Hfffffff4;
2571: data <= 32'Hfffffffb;
2572: data <= 32'Hfffffff3;
2573: data <= 32'Hfffffff7;
2574: data <= 32'Hfffffff8;
2575: data <= 32'Hfffffffa;
2576: data <= 32'Hfffffff6;
2577: data <= 32'Hfffffff6;
2578: data <= 32'Hfffffffb;
2579: data <= 32'Hfffffffa;
2580: data <= 32'Hfffffff9;
2581: data <= 32'Hfffffff2;
2582: data <= 32'Hffffffe9;
2583: data <= 32'Hffffffe6;
2584: data <= 32'Hfffffff6;
2585: data <= 32'Hfffffffc;
2586: data <= 32'Hfffffffa;
2587: data <= 32'Hfffffffc;
2588: data <= 32'Hfffffffc;
2589: data <= 32'Hfffffff9;
2590: data <= 32'H00000001;
2591: data <= 32'Hfffffff9;
2592: data <= 32'Hfffffff7;
2593: data <= 32'Hfffffff8;
2594: data <= 32'Hfffffff9;
2595: data <= 32'Hfffffffa;
2596: data <= 32'Hfffffff4;
2597: data <= 32'Hffffffef;
2598: data <= 32'Hffffffec;
2599: data <= 32'Hffffffe6;
2600: data <= 32'Hffffffe4;
2601: data <= 32'Hffffffe0;
2602: data <= 32'Hffffffe4;
2603: data <= 32'Hffffffe4;
2604: data <= 32'Hffffffea;
2605: data <= 32'Hffffffec;
2606: data <= 32'Hfffffff1;
2607: data <= 32'Hfffffff8;
2608: data <= 32'Hfffffff4;
2609: data <= 32'Hffffffe6;
2610: data <= 32'Hffffffd9;
2611: data <= 32'Hffffffdc;
2612: data <= 32'Hffffffe1;
2613: data <= 32'Hffffffe5;
2614: data <= 32'Hffffffe5;
2615: data <= 32'Hffffffe6;
2616: data <= 32'Hffffffdf;
2617: data <= 32'Hffffffde;
2618: data <= 32'Hffffffe6;
2619: data <= 32'Hffffffea;
2620: data <= 32'Hffffffeb;
2621: data <= 32'Hffffffec;
2622: data <= 32'Hffffffed;
2623: data <= 32'Hffffffec;
2624: data <= 32'Hfffffff1;
2625: data <= 32'Hfffffff2;
2626: data <= 32'Hfffffff4;
2627: data <= 32'Hfffffff5;
2628: data <= 32'Hfffffffa;
2629: data <= 32'Hfffffff8;
2630: data <= 32'Hfffffffa;
2631: data <= 32'Hfffffff5;
2632: data <= 32'Hffffffef;
2633: data <= 32'Hffffffef;
2634: data <= 32'Hffffffee;
2635: data <= 32'Hffffffef;
2636: data <= 32'Hfffffff0;
2637: data <= 32'Hffffffee;
2638: data <= 32'Hffffffec;
2639: data <= 32'Hffffffee;
2640: data <= 32'Hffffffec;
2641: data <= 32'Hffffffe7;
2642: data <= 32'Hffffffe9;
2643: data <= 32'Hffffffe3;
2644: data <= 32'Hffffffe2;
2645: data <= 32'Hffffffdb;
2646: data <= 32'Hffffffe2;
2647: data <= 32'Hffffffe0;
2648: data <= 32'Hffffffe6;
2649: data <= 32'Hffffffeb;
2650: data <= 32'Hfffffff0;
2651: data <= 32'Hffffffef;
2652: data <= 32'Hfffffff3;
2653: data <= 32'Hfffffff6;
2654: data <= 32'Hfffffff4;
2655: data <= 32'Hfffffff9;
2656: data <= 32'Hfffffff0;
2657: data <= 32'Hffffffef;
2658: data <= 32'Hffffffee;
2659: data <= 32'Hffffffe8;
2660: data <= 32'Hffffffe3;
2661: data <= 32'Hffffffea;
2662: data <= 32'Hffffffe9;
2663: data <= 32'Hfffffff5;
2664: data <= 32'Hfffffffb;
2665: data <= 32'Hfffffffb;
2666: data <= 32'Hfffffff9;
2667: data <= 32'Hfffffff3;
2668: data <= 32'Hfffffff6;
2669: data <= 32'H00000002;
2670: data <= 32'H00000007;
2671: data <= 32'H00000007;
2672: data <= 32'Hfffffffe;
2673: data <= 32'Hffffffeb;
2674: data <= 32'Hffffffdf;
2675: data <= 32'Hffffffd7;
2676: data <= 32'Hffffffdb;
2677: data <= 32'Hffffffe3;
2678: data <= 32'Hffffffec;
2679: data <= 32'Hffffffe7;
2680: data <= 32'Hffffffdb;
2681: data <= 32'Hffffffdd;
2682: data <= 32'Hffffffe8;
2683: data <= 32'Hfffffff5;
2684: data <= 32'H00000003;
2685: data <= 32'H0000000f;
2686: data <= 32'H00000012;
2687: data <= 32'H0000000d;
2688: data <= 32'H0000000a;
2689: data <= 32'H00000000;
2690: data <= 32'Hfffffffb;
2691: data <= 32'Hfffffffc;
2692: data <= 32'Hfffffffb;
2693: data <= 32'Hfffffffd;
2694: data <= 32'Hfffffffd;
2695: data <= 32'H00000000;
2696: data <= 32'H00000000;
2697: data <= 32'H00000001;
2698: data <= 32'H00000000;
2699: data <= 32'Hfffffffd;
2700: data <= 32'Hfffffffb;
2701: data <= 32'H00000001;
2702: data <= 32'Hffffffff;
2703: data <= 32'Hfffffffc;
2704: data <= 32'Hfffffffb;
2705: data <= 32'Hfffffffa;
2706: data <= 32'H00000000;
2707: data <= 32'Hfffffffd;
2708: data <= 32'Hfffffffd;
2709: data <= 32'Hfffffff9;
2710: data <= 32'Hfffffff4;
2711: data <= 32'Hfffffff4;
2712: data <= 32'H00000001;
2713: data <= 32'H00000006;
2714: data <= 32'H00000002;
2715: data <= 32'Hfffffffe;
2716: data <= 32'Hfffffffe;
2717: data <= 32'Hffffffff;
2718: data <= 32'Hffffffff;
2719: data <= 32'Hfffffffe;
2720: data <= 32'Hfffffff7;
2721: data <= 32'Hfffffff5;
2722: data <= 32'Hfffffff8;
2723: data <= 32'Hfffffff8;
2724: data <= 32'Hfffffff7;
2725: data <= 32'Hfffffff3;
2726: data <= 32'Hffffffef;
2727: data <= 32'Hffffffec;
2728: data <= 32'Hffffffe9;
2729: data <= 32'Hffffffe6;
2730: data <= 32'Hfffffff1;
2731: data <= 32'Hfffffff6;
2732: data <= 32'Hfffffff5;
2733: data <= 32'Hfffffffa;
2734: data <= 32'H00000000;
2735: data <= 32'Hfffffffe;
2736: data <= 32'Hfffffff0;
2737: data <= 32'Hffffffde;
2738: data <= 32'Hffffffd4;
2739: data <= 32'Hffffffda;
2740: data <= 32'Hffffffe4;
2741: data <= 32'Hffffffe3;
2742: data <= 32'Hffffffe5;
2743: data <= 32'Hffffffe4;
2744: data <= 32'Hffffffe6;
2745: data <= 32'Hffffffe8;
2746: data <= 32'Hfffffff2;
2747: data <= 32'Hfffffff1;
2748: data <= 32'Hffffffef;
2749: data <= 32'Hfffffff1;
2750: data <= 32'Hfffffff1;
2751: data <= 32'Hfffffff1;
2752: data <= 32'Hfffffff6;
2753: data <= 32'Hfffffffc;
2754: data <= 32'Hfffffffb;
2755: data <= 32'Hfffffff8;
2756: data <= 32'Hfffffffb;
2757: data <= 32'Hfffffff8;
2758: data <= 32'Hfffffff7;
2759: data <= 32'Hfffffff1;
2760: data <= 32'Hffffffef;
2761: data <= 32'Hffffffee;
2762: data <= 32'Hffffffed;
2763: data <= 32'Hfffffff2;
2764: data <= 32'Hffffffee;
2765: data <= 32'Hffffffed;
2766: data <= 32'Hfffffff1;
2767: data <= 32'Hfffffff2;
2768: data <= 32'Hfffffff2;
2769: data <= 32'Hffffffee;
2770: data <= 32'Hffffffeb;
2771: data <= 32'Hffffffe7;
2772: data <= 32'Hffffffe7;
2773: data <= 32'Hffffffe2;
2774: data <= 32'Hffffffe1;
2775: data <= 32'Hffffffe4;
2776: data <= 32'Hffffffe7;
2777: data <= 32'Hffffffe7;
2778: data <= 32'Hfffffff1;
2779: data <= 32'Hffffffef;
2780: data <= 32'Hffffffed;
2781: data <= 32'Hfffffff0;
2782: data <= 32'Hfffffff2;
2783: data <= 32'Hfffffff1;
2784: data <= 32'Hffffffef;
2785: data <= 32'Hffffffeb;
2786: data <= 32'Hffffffeb;
2787: data <= 32'Hffffffee;
2788: data <= 32'Hffffffe6;
2789: data <= 32'Hffffffe6;
2790: data <= 32'Hffffffe3;
2791: data <= 32'Hffffffea;
2792: data <= 32'Hfffffff6;
2793: data <= 32'Hfffffff8;
2794: data <= 32'Hfffffffa;
2795: data <= 32'Hfffffff6;
2796: data <= 32'Hffffffec;
2797: data <= 32'Hffffffef;
2798: data <= 32'Hfffffffe;
2799: data <= 32'Hfffffffe;
2800: data <= 32'Hfffffffb;
2801: data <= 32'Hfffffff7;
2802: data <= 32'Hffffffe6;
2803: data <= 32'Hffffffe6;
2804: data <= 32'Hffffffe7;
2805: data <= 32'Hffffffed;
2806: data <= 32'Hfffffff8;
2807: data <= 32'H00000002;
2808: data <= 32'Hfffffff7;
2809: data <= 32'Hfffffff8;
2810: data <= 32'Hfffffff2;
2811: data <= 32'Hfffffff6;
2812: data <= 32'H00000002;
2813: data <= 32'H00000007;
2814: data <= 32'H0000000d;
2815: data <= 32'H00000015;
2816: data <= 32'H00000013;
2817: data <= 32'Hfffffff5;
2818: data <= 32'Hfffffff2;
2819: data <= 32'Hfffffff4;
2820: data <= 32'Hfffffff1;
2821: data <= 32'Hfffffff2;
2822: data <= 32'Hfffffff5;
2823: data <= 32'Hfffffff5;
2824: data <= 32'Hfffffff4;
2825: data <= 32'Hfffffff1;
2826: data <= 32'Hfffffff5;
2827: data <= 32'Hfffffff1;
2828: data <= 32'Hfffffff2;
2829: data <= 32'Hfffffff3;
2830: data <= 32'Hfffffff5;
2831: data <= 32'Hffffffec;
2832: data <= 32'Hfffffff0;
2833: data <= 32'Hfffffff0;
2834: data <= 32'Hffffffee;
2835: data <= 32'Hffffffe9;
2836: data <= 32'Hffffffe6;
2837: data <= 32'Hffffffe2;
2838: data <= 32'Hffffffe6;
2839: data <= 32'Hffffffeb;
2840: data <= 32'Hfffffff0;
2841: data <= 32'Hfffffff2;
2842: data <= 32'Hffffffec;
2843: data <= 32'Hffffffea;
2844: data <= 32'Hffffffed;
2845: data <= 32'Hfffffff2;
2846: data <= 32'Hffffffef;
2847: data <= 32'Hfffffff5;
2848: data <= 32'Hfffffff1;
2849: data <= 32'Hfffffff2;
2850: data <= 32'Hfffffff3;
2851: data <= 32'Hfffffff6;
2852: data <= 32'Hfffffff4;
2853: data <= 32'Hfffffff3;
2854: data <= 32'Hffffffeb;
2855: data <= 32'Hffffffe5;
2856: data <= 32'Hffffffe4;
2857: data <= 32'Hffffffec;
2858: data <= 32'Hfffffff5;
2859: data <= 32'Hfffffffb;
2860: data <= 32'Hfffffffb;
2861: data <= 32'H00000001;
2862: data <= 32'H00000003;
2863: data <= 32'Hfffffffa;
2864: data <= 32'Hffffffe6;
2865: data <= 32'Hffffffd5;
2866: data <= 32'Hffffffd1;
2867: data <= 32'Hffffffd4;
2868: data <= 32'Hffffffda;
2869: data <= 32'Hffffffda;
2870: data <= 32'Hffffffdc;
2871: data <= 32'Hffffffd9;
2872: data <= 32'Hffffffea;
2873: data <= 32'Hffffffeb;
2874: data <= 32'Hffffffec;
2875: data <= 32'Hffffffeb;
2876: data <= 32'Hffffffe6;
2877: data <= 32'Hffffffe3;
2878: data <= 32'Hffffffe7;
2879: data <= 32'Hffffffea;
2880: data <= 32'Hffffffec;
2881: data <= 32'Hfffffff1;
2882: data <= 32'Hfffffff2;
2883: data <= 32'Hffffffee;
2884: data <= 32'Hfffffff1;
2885: data <= 32'Hffffffed;
2886: data <= 32'Hffffffec;
2887: data <= 32'Hffffffea;
2888: data <= 32'Hffffffe7;
2889: data <= 32'Hffffffe8;
2890: data <= 32'Hffffffeb;
2891: data <= 32'Hffffffe7;
2892: data <= 32'Hffffffe6;
2893: data <= 32'Hffffffe9;
2894: data <= 32'Hffffffe8;
2895: data <= 32'Hffffffe7;
2896: data <= 32'Hffffffe9;
2897: data <= 32'Hffffffe6;
2898: data <= 32'Hffffffe2;
2899: data <= 32'Hffffffe0;
2900: data <= 32'Hffffffde;
2901: data <= 32'Hffffffdd;
2902: data <= 32'Hffffffda;
2903: data <= 32'Hffffffdd;
2904: data <= 32'Hffffffd5;
2905: data <= 32'Hffffffd9;
2906: data <= 32'Hffffffda;
2907: data <= 32'Hffffffdf;
2908: data <= 32'Hffffffe0;
2909: data <= 32'Hffffffdf;
2910: data <= 32'Hffffffe0;
2911: data <= 32'Hffffffde;
2912: data <= 32'Hffffffdd;
2913: data <= 32'Hffffffdb;
2914: data <= 32'Hffffffdb;
2915: data <= 32'Hffffffdd;
2916: data <= 32'Hffffffdf;
2917: data <= 32'Hffffffdd;
2918: data <= 32'Hffffffe0;
2919: data <= 32'Hffffffe4;
2920: data <= 32'Hffffffe8;
2921: data <= 32'Hfffffff3;
2922: data <= 32'Hfffffffc;
2923: data <= 32'Hfffffff6;
2924: data <= 32'Hffffffee;
2925: data <= 32'Hffffffee;
2926: data <= 32'Hffffffeb;
2927: data <= 32'Hfffffff7;
2928: data <= 32'Hfffffff8;
2929: data <= 32'Hfffffffb;
2930: data <= 32'Hfffffffe;
2931: data <= 32'Hfffffff9;
2932: data <= 32'Hfffffff8;
2933: data <= 32'Hfffffffe;
2934: data <= 32'Hfffffffe;
2935: data <= 32'H00000004;
2936: data <= 32'H00000005;
2937: data <= 32'Hfffffffd;
2938: data <= 32'Hfffffff8;
2939: data <= 32'Hfffffff4;
2940: data <= 32'Hfffffff6;
2941: data <= 32'Hfffffff4;
2942: data <= 32'Hfffffffb;
2943: data <= 32'Hfffffffe;
2944: data <= 32'H0000000b;
2945: data <= 32'Hfffffffe;
2946: data <= 32'Hfffffffb;
2947: data <= 32'Hfffffff7;
2948: data <= 32'Hfffffff8;
2949: data <= 32'Hfffffff5;
2950: data <= 32'Hfffffff6;
2951: data <= 32'Hfffffff4;
2952: data <= 32'Hfffffff5;
2953: data <= 32'Hfffffff4;
2954: data <= 32'Hfffffff4;
2955: data <= 32'Hfffffff5;
2956: data <= 32'Hfffffffb;
2957: data <= 32'Hfffffff5;
2958: data <= 32'Hfffffff2;
2959: data <= 32'Hfffffff4;
2960: data <= 32'Hffffffeb;
2961: data <= 32'Hffffffe8;
2962: data <= 32'Hffffffec;
2963: data <= 32'Hffffffe5;
2964: data <= 32'Hffffffe5;
2965: data <= 32'Hffffffe6;
2966: data <= 32'Hffffffea;
2967: data <= 32'Hfffffff4;
2968: data <= 32'Hfffffff5;
2969: data <= 32'Hfffffff4;
2970: data <= 32'Hffffffee;
2971: data <= 32'Hfffffff1;
2972: data <= 32'Hfffffff3;
2973: data <= 32'Hfffffff6;
2974: data <= 32'Hfffffffa;
2975: data <= 32'Hfffffffd;
2976: data <= 32'Hfffffffb;
2977: data <= 32'Hfffffffc;
2978: data <= 32'Hfffffffd;
2979: data <= 32'Hfffffffd;
2980: data <= 32'Hfffffffc;
2981: data <= 32'Hfffffff9;
2982: data <= 32'Hffffffee;
2983: data <= 32'Hffffffe7;
2984: data <= 32'Hffffffea;
2985: data <= 32'Hfffffff1;
2986: data <= 32'Hfffffff6;
2987: data <= 32'Hfffffffb;
2988: data <= 32'H00000002;
2989: data <= 32'H00000002;
2990: data <= 32'Hfffffffb;
2991: data <= 32'Hffffffee;
2992: data <= 32'Hffffffdd;
2993: data <= 32'Hffffffd5;
2994: data <= 32'Hffffffd7;
2995: data <= 32'Hffffffdb;
2996: data <= 32'Hffffffde;
2997: data <= 32'Hffffffd8;
2998: data <= 32'Hffffffde;
2999: data <= 32'Hffffffe0;
3000: data <= 32'Hffffffea;
3001: data <= 32'Hffffffeb;
3002: data <= 32'Hffffffed;
3003: data <= 32'Hffffffe8;
3004: data <= 32'Hffffffe4;
3005: data <= 32'Hffffffe7;
3006: data <= 32'Hffffffe8;
3007: data <= 32'Hffffffec;
3008: data <= 32'Hfffffff1;
3009: data <= 32'Hffffffee;
3010: data <= 32'Hffffffed;
3011: data <= 32'Hfffffff0;
3012: data <= 32'Hffffffeb;
3013: data <= 32'Hffffffe9;
3014: data <= 32'Hffffffec;
3015: data <= 32'Hffffffe4;
3016: data <= 32'Hffffffe7;
3017: data <= 32'Hffffffe7;
3018: data <= 32'Hffffffe6;
3019: data <= 32'Hffffffe5;
3020: data <= 32'Hffffffec;
3021: data <= 32'Hffffffec;
3022: data <= 32'Hffffffed;
3023: data <= 32'Hfffffff1;
3024: data <= 32'Hffffffef;
3025: data <= 32'Hffffffeb;
3026: data <= 32'Hffffffe7;
3027: data <= 32'Hffffffe5;
3028: data <= 32'Hffffffe0;
3029: data <= 32'Hffffffe5;
3030: data <= 32'Hffffffe0;
3031: data <= 32'Hffffffe0;
3032: data <= 32'Hffffffe2;
3033: data <= 32'Hffffffe1;
3034: data <= 32'Hffffffe1;
3035: data <= 32'Hffffffe6;
3036: data <= 32'Hffffffe7;
3037: data <= 32'Hffffffe5;
3038: data <= 32'Hffffffe3;
3039: data <= 32'Hffffffe3;
3040: data <= 32'Hffffffe2;
3041: data <= 32'Hffffffdf;
3042: data <= 32'Hffffffe1;
3043: data <= 32'Hffffffe5;
3044: data <= 32'Hffffffe6;
3045: data <= 32'Hffffffe6;
3046: data <= 32'Hffffffec;
3047: data <= 32'Hffffffe9;
3048: data <= 32'Hffffffeb;
3049: data <= 32'Hfffffff4;
3050: data <= 32'Hfffffff7;
3051: data <= 32'Hfffffffc;
3052: data <= 32'Hfffffff8;
3053: data <= 32'Hfffffff5;
3054: data <= 32'Hfffffff2;
3055: data <= 32'Hfffffff3;
3056: data <= 32'Hfffffff5;
3057: data <= 32'H00000002;
3058: data <= 32'H00000005;
3059: data <= 32'H00000005;
3060: data <= 32'H00000009;
3061: data <= 32'H00000007;
3062: data <= 32'H00000007;
3063: data <= 32'Hffffffff;
3064: data <= 32'Hfffffffe;
3065: data <= 32'H00000000;
3066: data <= 32'H00000000;
3067: data <= 32'Hfffffff1;
3068: data <= 32'Hfffffff4;
3069: data <= 32'Hfffffff4;
3070: data <= 32'Hfffffff3;
3071: data <= 32'Hfffffffa;
3072: data <= 32'H00000000;
3073: data <= 32'H00000000;
3074: data <= 32'H00000002;
3075: data <= 32'Hfffffffc;
3076: data <= 32'Hfffffffd;
3077: data <= 32'Hfffffffa;
3078: data <= 32'Hfffffff9;
3079: data <= 32'Hfffffff6;
3080: data <= 32'Hfffffff8;
3081: data <= 32'Hfffffffa;
3082: data <= 32'Hfffffffd;
3083: data <= 32'H00000004;
3084: data <= 32'H00000007;
3085: data <= 32'H00000005;
3086: data <= 32'H00000004;
3087: data <= 32'Hfffffffc;
3088: data <= 32'Hfffffff3;
3089: data <= 32'Hfffffff1;
3090: data <= 32'Hffffffef;
3091: data <= 32'Hfffffff0;
3092: data <= 32'Hfffffff7;
3093: data <= 32'Hfffffff5;
3094: data <= 32'Hfffffffc;
3095: data <= 32'H00000000;
3096: data <= 32'H00000002;
3097: data <= 32'Hfffffffe;
3098: data <= 32'Hfffffffa;
3099: data <= 32'Hfffffffc;
3100: data <= 32'Hfffffffb;
3101: data <= 32'Hfffffffd;
3102: data <= 32'Hffffffff;
3103: data <= 32'Hfffffffe;
3104: data <= 32'Hfffffffc;
3105: data <= 32'Hfffffffb;
3106: data <= 32'Hfffffff9;
3107: data <= 32'Hffffffff;
3108: data <= 32'Hfffffff8;
3109: data <= 32'Hfffffff1;
3110: data <= 32'Hffffffe8;
3111: data <= 32'Hffffffea;
3112: data <= 32'Hffffffec;
3113: data <= 32'Hfffffff1;
3114: data <= 32'Hfffffff8;
3115: data <= 32'Hfffffffd;
3116: data <= 32'H00000003;
3117: data <= 32'H00000003;
3118: data <= 32'Hfffffff5;
3119: data <= 32'Hffffffe5;
3120: data <= 32'Hffffffe3;
3121: data <= 32'Hffffffe2;
3122: data <= 32'Hffffffea;
3123: data <= 32'Hffffffee;
3124: data <= 32'Hffffffeb;
3125: data <= 32'Hffffffe9;
3126: data <= 32'Hfffffff0;
3127: data <= 32'Hfffffff1;
3128: data <= 32'Hfffffff4;
3129: data <= 32'Hfffffff4;
3130: data <= 32'Hffffffef;
3131: data <= 32'Hfffffff0;
3132: data <= 32'Hffffffef;
3133: data <= 32'Hfffffff0;
3134: data <= 32'Hfffffff5;
3135: data <= 32'Hfffffff2;
3136: data <= 32'Hfffffff6;
3137: data <= 32'Hfffffff5;
3138: data <= 32'Hfffffff0;
3139: data <= 32'Hfffffff0;
3140: data <= 32'Hfffffff6;
3141: data <= 32'Hfffffff0;
3142: data <= 32'Hffffffec;
3143: data <= 32'Hffffffeb;
3144: data <= 32'Hffffffec;
3145: data <= 32'Hffffffe6;
3146: data <= 32'Hffffffe9;
3147: data <= 32'Hffffffe7;
3148: data <= 32'Hffffffea;
3149: data <= 32'Hfffffff4;
3150: data <= 32'Hfffffff6;
3151: data <= 32'Hfffffff9;
3152: data <= 32'Hfffffffa;
3153: data <= 32'Hfffffff8;
3154: data <= 32'Hfffffff4;
3155: data <= 32'Hfffffff1;
3156: data <= 32'Hffffffeb;
3157: data <= 32'Hffffffe8;
3158: data <= 32'Hffffffe7;
3159: data <= 32'Hffffffe7;
3160: data <= 32'Hffffffe8;
3161: data <= 32'Hffffffe9;
3162: data <= 32'Hffffffec;
3163: data <= 32'Hfffffff0;
3164: data <= 32'Hfffffff2;
3165: data <= 32'Hfffffff3;
3166: data <= 32'Hfffffff6;
3167: data <= 32'Hfffffff5;
3168: data <= 32'Hffffffef;
3169: data <= 32'Hfffffff2;
3170: data <= 32'Hffffffee;
3171: data <= 32'Hffffffed;
3172: data <= 32'Hffffffef;
3173: data <= 32'Hffffffed;
3174: data <= 32'Hffffffec;
3175: data <= 32'Hffffffeb;
3176: data <= 32'Hffffffe5;
3177: data <= 32'Hffffffe1;
3178: data <= 32'Hffffffe6;
3179: data <= 32'Hffffffeb;
3180: data <= 32'Hffffffea;
3181: data <= 32'Hffffffeb;
3182: data <= 32'Hffffffe6;
3183: data <= 32'Hffffffe0;
3184: data <= 32'Hffffffe3;
3185: data <= 32'Hffffffed;
3186: data <= 32'Hfffffff5;
3187: data <= 32'Hfffffffa;
3188: data <= 32'Hfffffffc;
3189: data <= 32'Hfffffffd;
3190: data <= 32'H00000001;
3191: data <= 32'Hfffffff7;
3192: data <= 32'Hfffffff0;
3193: data <= 32'Hfffffff3;
3194: data <= 32'Hfffffff8;
3195: data <= 32'Hfffffff5;
3196: data <= 32'Hffffffec;
3197: data <= 32'Hfffffff4;
3198: data <= 32'Hfffffff7;
3199: data <= 32'Hfffffffb;
3200: data <= 32'Hfffffffc;
3201: data <= 32'H00000003;
3202: data <= 32'H00000006;
3203: data <= 32'H00000003;
3204: data <= 32'Hffffffff;
3205: data <= 32'H00000000;
3206: data <= 32'H00000001;
3207: data <= 32'Hfffffffc;
3208: data <= 32'H00000003;
3209: data <= 32'H00000007;
3210: data <= 32'H00000010;
3211: data <= 32'H00000013;
3212: data <= 32'H00000017;
3213: data <= 32'H0000001a;
3214: data <= 32'H00000014;
3215: data <= 32'H0000000c;
3216: data <= 32'H00000004;
3217: data <= 32'H00000002;
3218: data <= 32'H00000004;
3219: data <= 32'H00000004;
3220: data <= 32'H00000007;
3221: data <= 32'H00000009;
3222: data <= 32'H0000000d;
3223: data <= 32'H0000000c;
3224: data <= 32'H0000000c;
3225: data <= 32'H00000006;
3226: data <= 32'H00000002;
3227: data <= 32'H00000001;
3228: data <= 32'H00000002;
3229: data <= 32'H00000000;
3230: data <= 32'H00000000;
3231: data <= 32'Hffffffff;
3232: data <= 32'Hfffffffb;
3233: data <= 32'Hfffffffd;
3234: data <= 32'H00000002;
3235: data <= 32'H00000004;
3236: data <= 32'Hfffffff9;
3237: data <= 32'Hfffffff2;
3238: data <= 32'Hffffffef;
3239: data <= 32'Hfffffff5;
3240: data <= 32'Hfffffffa;
3241: data <= 32'Hfffffffe;
3242: data <= 32'Hffffffff;
3243: data <= 32'H00000005;
3244: data <= 32'H0000000c;
3245: data <= 32'Hffffffff;
3246: data <= 32'Hfffffff0;
3247: data <= 32'Hffffffe2;
3248: data <= 32'Hffffffe6;
3249: data <= 32'Hffffffea;
3250: data <= 32'Hffffffef;
3251: data <= 32'Hffffffef;
3252: data <= 32'Hfffffff0;
3253: data <= 32'Hfffffff2;
3254: data <= 32'Hfffffff6;
3255: data <= 32'Hfffffffc;
3256: data <= 32'Hfffffff9;
3257: data <= 32'Hfffffff8;
3258: data <= 32'Hfffffff3;
3259: data <= 32'Hfffffff2;
3260: data <= 32'Hfffffff3;
3261: data <= 32'Hfffffff6;
3262: data <= 32'Hfffffff4;
3263: data <= 32'Hfffffff5;
3264: data <= 32'Hfffffffb;
3265: data <= 32'Hfffffff7;
3266: data <= 32'Hfffffff7;
3267: data <= 32'Hfffffffa;
3268: data <= 32'Hfffffff6;
3269: data <= 32'Hfffffff6;
3270: data <= 32'Hfffffff5;
3271: data <= 32'Hfffffff1;
3272: data <= 32'Hfffffff1;
3273: data <= 32'Hffffffee;
3274: data <= 32'Hffffffec;
3275: data <= 32'Hffffffec;
3276: data <= 32'Hffffffef;
3277: data <= 32'Hfffffff5;
3278: data <= 32'Hfffffff8;
3279: data <= 32'Hfffffffb;
3280: data <= 32'Hfffffffc;
3281: data <= 32'Hfffffffe;
3282: data <= 32'Hfffffffa;
3283: data <= 32'Hfffffff5;
3284: data <= 32'Hfffffff0;
3285: data <= 32'Hffffffea;
3286: data <= 32'Hffffffeb;
3287: data <= 32'Hffffffeb;
3288: data <= 32'Hffffffe9;
3289: data <= 32'Hffffffec;
3290: data <= 32'Hfffffff2;
3291: data <= 32'Hfffffff4;
3292: data <= 32'Hfffffff8;
3293: data <= 32'Hfffffffe;
3294: data <= 32'Hfffffffd;
3295: data <= 32'Hfffffffe;
3296: data <= 32'Hfffffffd;
3297: data <= 32'Hfffffffd;
3298: data <= 32'Hfffffff8;
3299: data <= 32'Hfffffff9;
3300: data <= 32'Hfffffff8;
3301: data <= 32'Hfffffff5;
3302: data <= 32'Hfffffff1;
3303: data <= 32'Hffffffee;
3304: data <= 32'Hffffffe6;
3305: data <= 32'Hffffffe0;
3306: data <= 32'Hffffffdf;
3307: data <= 32'Hffffffe1;
3308: data <= 32'Hffffffe7;
3309: data <= 32'Hffffffe8;
3310: data <= 32'Hffffffe3;
3311: data <= 32'Hffffffe0;
3312: data <= 32'Hffffffe1;
3313: data <= 32'Hffffffe7;
3314: data <= 32'Hfffffff3;
3315: data <= 32'Hfffffffb;
3316: data <= 32'Hfffffffd;
3317: data <= 32'H00000000;
3318: data <= 32'H00000004;
3319: data <= 32'H00000004;
3320: data <= 32'Hfffffffc;
3321: data <= 32'Hfffffff7;
3322: data <= 32'Hffffffff;
3323: data <= 32'H00000006;
3324: data <= 32'Hfffffffc;
3325: data <= 32'Hfffffffd;
3326: data <= 32'Hfffffffb;
3327: data <= 32'H00000001;
3328: data <= 32'H00000005;
3329: data <= 32'H00000005;
3330: data <= 32'Hffffffff;
3331: data <= 32'H00000000;
3332: data <= 32'Hfffffffc;
3333: data <= 32'Hfffffffd;
3334: data <= 32'Hffffffff;
3335: data <= 32'Hffffffff;
3336: data <= 32'H00000001;
3337: data <= 32'H0000000d;
3338: data <= 32'H00000013;
3339: data <= 32'H00000015;
3340: data <= 32'H0000001a;
3341: data <= 32'H00000017;
3342: data <= 32'H00000013;
3343: data <= 32'H00000008;
3344: data <= 32'H00000001;
3345: data <= 32'H00000005;
3346: data <= 32'H00000007;
3347: data <= 32'H00000006;
3348: data <= 32'H00000006;
3349: data <= 32'H00000009;
3350: data <= 32'H0000000b;
3351: data <= 32'H00000008;
3352: data <= 32'H00000007;
3353: data <= 32'H00000004;
3354: data <= 32'H00000004;
3355: data <= 32'H00000003;
3356: data <= 32'H00000002;
3357: data <= 32'H00000006;
3358: data <= 32'H00000002;
3359: data <= 32'H00000000;
3360: data <= 32'H00000001;
3361: data <= 32'H0000000b;
3362: data <= 32'H00000010;
3363: data <= 32'H00000010;
3364: data <= 32'H00000003;
3365: data <= 32'Hfffffffc;
3366: data <= 32'Hffffffff;
3367: data <= 32'H00000008;
3368: data <= 32'H00000011;
3369: data <= 32'H0000000d;
3370: data <= 32'H0000000a;
3371: data <= 32'H00000013;
3372: data <= 32'H00000012;
3373: data <= 32'Hffffffff;
3374: data <= 32'Hfffffff0;
3375: data <= 32'Hffffffe2;
3376: data <= 32'Hffffffe7;
3377: data <= 32'Hffffffe9;
3378: data <= 32'Hffffffee;
3379: data <= 32'Hfffffff0;
3380: data <= 32'Hffffffef;
3381: data <= 32'Hfffffff4;
3382: data <= 32'Hfffffff7;
3383: data <= 32'Hfffffff6;
3384: data <= 32'Hfffffff5;
3385: data <= 32'Hfffffff4;
3386: data <= 32'Hffffffed;
3387: data <= 32'Hfffffff0;
3388: data <= 32'Hfffffff2;
3389: data <= 32'Hfffffff0;
3390: data <= 32'Hfffffff1;
3391: data <= 32'Hfffffff4;
3392: data <= 32'Hfffffff3;
3393: data <= 32'Hfffffff6;
3394: data <= 32'Hfffffff7;
3395: data <= 32'Hfffffff5;
3396: data <= 32'Hfffffff6;
3397: data <= 32'Hfffffff7;
3398: data <= 32'Hfffffff5;
3399: data <= 32'Hfffffff3;
3400: data <= 32'Hfffffff5;
3401: data <= 32'Hfffffff1;
3402: data <= 32'Hfffffff2;
3403: data <= 32'Hfffffff1;
3404: data <= 32'Hfffffff4;
3405: data <= 32'Hfffffff8;
3406: data <= 32'Hfffffff8;
3407: data <= 32'Hfffffffa;
3408: data <= 32'Hfffffffb;
3409: data <= 32'Hfffffff9;
3410: data <= 32'Hfffffffa;
3411: data <= 32'Hfffffff6;
3412: data <= 32'Hfffffff2;
3413: data <= 32'Hffffffef;
3414: data <= 32'Hfffffff1;
3415: data <= 32'Hffffffee;
3416: data <= 32'Hfffffff0;
3417: data <= 32'Hfffffff2;
3418: data <= 32'Hfffffff4;
3419: data <= 32'Hfffffff8;
3420: data <= 32'Hfffffffd;
3421: data <= 32'Hfffffffd;
3422: data <= 32'Hfffffffd;
3423: data <= 32'H00000002;
3424: data <= 32'H00000002;
3425: data <= 32'H00000001;
3426: data <= 32'H00000001;
3427: data <= 32'H00000000;
3428: data <= 32'Hfffffffc;
3429: data <= 32'Hfffffffc;
3430: data <= 32'Hfffffff7;
3431: data <= 32'Hffffffed;
3432: data <= 32'Hffffffe9;
3433: data <= 32'Hffffffe3;
3434: data <= 32'Hffffffd9;
3435: data <= 32'Hffffffdf;
3436: data <= 32'Hffffffe4;
3437: data <= 32'Hffffffe7;
3438: data <= 32'Hffffffeb;
3439: data <= 32'Hffffffe7;
3440: data <= 32'Hffffffe8;
3441: data <= 32'Hfffffff2;
3442: data <= 32'Hfffffffb;
3443: data <= 32'H00000006;
3444: data <= 32'H00000009;
3445: data <= 32'H00000008;
3446: data <= 32'H00000008;
3447: data <= 32'H0000000f;
3448: data <= 32'H00000009;
3449: data <= 32'H00000005;
3450: data <= 32'H0000000a;
3451: data <= 32'H00000012;
3452: data <= 32'H00000011;
3453: data <= 32'H00000005;
3454: data <= 32'H00000002;
3455: data <= 32'H00000005;
3456: data <= 32'H00000005;
3457: data <= 32'H00000002;
3458: data <= 32'H00000000;
3459: data <= 32'Hffffffff;
3460: data <= 32'Hfffffffe;
3461: data <= 32'Hffffffff;
3462: data <= 32'Hfffffffe;
3463: data <= 32'H00000002;
3464: data <= 32'H00000003;
3465: data <= 32'H00000008;
3466: data <= 32'H00000014;
3467: data <= 32'H00000016;
3468: data <= 32'H00000016;
3469: data <= 32'H00000016;
3470: data <= 32'H0000000b;
3471: data <= 32'Hffffffff;
3472: data <= 32'Hfffffffb;
3473: data <= 32'H00000000;
3474: data <= 32'H00000005;
3475: data <= 32'H00000004;
3476: data <= 32'H00000003;
3477: data <= 32'H00000003;
3478: data <= 32'H00000003;
3479: data <= 32'Hffffffff;
3480: data <= 32'Hffffffff;
3481: data <= 32'H00000000;
3482: data <= 32'H00000002;
3483: data <= 32'H00000004;
3484: data <= 32'H00000006;
3485: data <= 32'H00000004;
3486: data <= 32'H00000000;
3487: data <= 32'Hfffffffb;
3488: data <= 32'Hfffffffd;
3489: data <= 32'H00000009;
3490: data <= 32'H0000000b;
3491: data <= 32'H00000005;
3492: data <= 32'Hfffffffd;
3493: data <= 32'Hfffffff9;
3494: data <= 32'Hfffffffc;
3495: data <= 32'H00000007;
3496: data <= 32'H0000000a;
3497: data <= 32'H00000008;
3498: data <= 32'H0000000b;
3499: data <= 32'H0000000f;
3500: data <= 32'H0000000f;
3501: data <= 32'Hfffffffd;
3502: data <= 32'Hffffffef;
3503: data <= 32'Hffffffea;
3504: data <= 32'Hffffffea;
3505: data <= 32'Hffffffef;
3506: data <= 32'Hfffffff5;
3507: data <= 32'Hfffffff5;
3508: data <= 32'Hfffffff8;
3509: data <= 32'Hfffffffc;
3510: data <= 32'Hffffffff;
3511: data <= 32'H00000001;
3512: data <= 32'Hfffffff9;
3513: data <= 32'Hfffffff6;
3514: data <= 32'Hfffffff7;
3515: data <= 32'Hfffffff5;
3516: data <= 32'Hfffffff6;
3517: data <= 32'Hfffffff7;
3518: data <= 32'Hfffffff6;
3519: data <= 32'Hfffffff6;
3520: data <= 32'Hfffffff5;
3521: data <= 32'Hfffffff3;
3522: data <= 32'Hfffffff5;
3523: data <= 32'Hfffffff4;
3524: data <= 32'Hfffffff2;
3525: data <= 32'Hfffffff5;
3526: data <= 32'Hfffffff2;
3527: data <= 32'Hfffffff1;
3528: data <= 32'Hfffffff2;
3529: data <= 32'Hfffffff2;
3530: data <= 32'Hfffffff4;
3531: data <= 32'Hfffffff1;
3532: data <= 32'Hffffffef;
3533: data <= 32'Hffffffee;
3534: data <= 32'Hfffffff1;
3535: data <= 32'Hffffffee;
3536: data <= 32'Hffffffef;
3537: data <= 32'Hffffffee;
3538: data <= 32'Hffffffeb;
3539: data <= 32'Hffffffea;
3540: data <= 32'Hffffffe9;
3541: data <= 32'Hffffffea;
3542: data <= 32'Hffffffe8;
3543: data <= 32'Hffffffe9;
3544: data <= 32'Hffffffed;
3545: data <= 32'Hffffffed;
3546: data <= 32'Hfffffff1;
3547: data <= 32'Hfffffff5;
3548: data <= 32'Hfffffff7;
3549: data <= 32'Hfffffff8;
3550: data <= 32'Hfffffff7;
3551: data <= 32'Hfffffff9;
3552: data <= 32'Hfffffffc;
3553: data <= 32'Hfffffffd;
3554: data <= 32'Hffffffff;
3555: data <= 32'Hffffffff;
3556: data <= 32'Hfffffffe;
3557: data <= 32'Hfffffffb;
3558: data <= 32'Hfffffff8;
3559: data <= 32'Hfffffff3;
3560: data <= 32'Hffffffef;
3561: data <= 32'Hffffffed;
3562: data <= 32'Hffffffe9;
3563: data <= 32'Hffffffe6;
3564: data <= 32'Hffffffeb;
3565: data <= 32'Hfffffff3;
3566: data <= 32'Hfffffff2;
3567: data <= 32'Hfffffff3;
3568: data <= 32'Hfffffff5;
3569: data <= 32'Hfffffffd;
3570: data <= 32'H00000006;
3571: data <= 32'H0000000d;
3572: data <= 32'H00000012;
3573: data <= 32'H00000013;
3574: data <= 32'H00000008;
3575: data <= 32'H00000009;
3576: data <= 32'H0000000a;
3577: data <= 32'H00000002;
3578: data <= 32'H00000005;
3579: data <= 32'H00000010;
3580: data <= 32'H0000000c;
3581: data <= 32'H00000007;
3582: data <= 32'H00000002;
3583: data <= 32'Hfffffff9;
3584: data <= 32'Hfffffffc;
3585: data <= 32'H00000005;
3586: data <= 32'H00000000;
3587: data <= 32'H00000001;
3588: data <= 32'H00000001;
3589: data <= 32'Hfffffffd;
3590: data <= 32'Hffffffff;
3591: data <= 32'H00000001;
3592: data <= 32'H00000001;
3593: data <= 32'H0000000a;
3594: data <= 32'H00000011;
3595: data <= 32'H00000014;
3596: data <= 32'H0000001a;
3597: data <= 32'H00000011;
3598: data <= 32'H00000009;
3599: data <= 32'H00000002;
3600: data <= 32'H00000001;
3601: data <= 32'H00000005;
3602: data <= 32'H00000008;
3603: data <= 32'H0000000b;
3604: data <= 32'H00000007;
3605: data <= 32'H00000006;
3606: data <= 32'H00000006;
3607: data <= 32'H00000002;
3608: data <= 32'H00000000;
3609: data <= 32'H00000002;
3610: data <= 32'H00000004;
3611: data <= 32'H00000001;
3612: data <= 32'H00000001;
3613: data <= 32'H00000001;
3614: data <= 32'Hfffffffa;
3615: data <= 32'Hfffffff2;
3616: data <= 32'Hfffffff6;
3617: data <= 32'Hfffffffd;
3618: data <= 32'H00000002;
3619: data <= 32'Hfffffff6;
3620: data <= 32'Hfffffff2;
3621: data <= 32'Hfffffff1;
3622: data <= 32'Hfffffff4;
3623: data <= 32'Hfffffffa;
3624: data <= 32'Hfffffffc;
3625: data <= 32'Hfffffffd;
3626: data <= 32'Hfffffffe;
3627: data <= 32'H00000001;
3628: data <= 32'H00000002;
3629: data <= 32'Hfffffff9;
3630: data <= 32'Hfffffff1;
3631: data <= 32'Hffffffec;
3632: data <= 32'Hfffffff1;
3633: data <= 32'Hfffffff4;
3634: data <= 32'Hfffffff7;
3635: data <= 32'Hfffffff9;
3636: data <= 32'Hffffffff;
3637: data <= 32'H00000006;
3638: data <= 32'H0000000a;
3639: data <= 32'H00000007;
3640: data <= 32'H00000006;
3641: data <= 32'H00000001;
3642: data <= 32'H00000000;
3643: data <= 32'Hfffffffd;
3644: data <= 32'H00000000;
3645: data <= 32'Hfffffffd;
3646: data <= 32'Hfffffffe;
3647: data <= 32'Hfffffffd;
3648: data <= 32'Hfffffffb;
3649: data <= 32'Hfffffffa;
3650: data <= 32'Hfffffff9;
3651: data <= 32'Hfffffff8;
3652: data <= 32'Hfffffff6;
3653: data <= 32'Hfffffff5;
3654: data <= 32'Hfffffff6;
3655: data <= 32'Hfffffff3;
3656: data <= 32'Hfffffff5;
3657: data <= 32'Hfffffff5;
3658: data <= 32'Hfffffff7;
3659: data <= 32'Hfffffff6;
3660: data <= 32'Hfffffff6;
3661: data <= 32'Hfffffff1;
3662: data <= 32'Hfffffff3;
3663: data <= 32'Hfffffff0;
3664: data <= 32'Hffffffef;
3665: data <= 32'Hffffffee;
3666: data <= 32'Hffffffea;
3667: data <= 32'Hffffffe9;
3668: data <= 32'Hffffffe8;
3669: data <= 32'Hffffffeb;
3670: data <= 32'Hffffffea;
3671: data <= 32'Hffffffec;
3672: data <= 32'Hffffffef;
3673: data <= 32'Hfffffff1;
3674: data <= 32'Hfffffff1;
3675: data <= 32'Hfffffff3;
3676: data <= 32'Hfffffff5;
3677: data <= 32'Hfffffff5;
3678: data <= 32'Hfffffff3;
3679: data <= 32'Hfffffff4;
3680: data <= 32'Hfffffff7;
3681: data <= 32'Hfffffff7;
3682: data <= 32'Hfffffff6;
3683: data <= 32'Hfffffff9;
3684: data <= 32'Hfffffff9;
3685: data <= 32'Hfffffff9;
3686: data <= 32'Hfffffff8;
3687: data <= 32'Hfffffff2;
3688: data <= 32'Hfffffff0;
3689: data <= 32'Hfffffff6;
3690: data <= 32'Hfffffff0;
3691: data <= 32'Hfffffff1;
3692: data <= 32'Hfffffff3;
3693: data <= 32'Hfffffff9;
3694: data <= 32'Hfffffffb;
3695: data <= 32'Hfffffff6;
3696: data <= 32'Hfffffff8;
3697: data <= 32'H00000004;
3698: data <= 32'H0000000a;
3699: data <= 32'H00000011;
3700: data <= 32'H00000015;
3701: data <= 32'H00000011;
3702: data <= 32'H0000000a;
3703: data <= 32'H00000004;
3704: data <= 32'H00000001;
3705: data <= 32'H00000001;
3706: data <= 32'Hfffffffe;
3707: data <= 32'H00000006;
3708: data <= 32'H0000000a;
3709: data <= 32'H00000004;
3710: data <= 32'Hfffffffb;
3711: data <= 32'Hfffffff6;
3712: data <= 32'Hffffffea;
3713: data <= 32'Hfffffffa;
3714: data <= 32'Hfffffffc;
3715: data <= 32'Hfffffffa;
3716: data <= 32'Hfffffff9;
3717: data <= 32'Hfffffffa;
3718: data <= 32'Hfffffff5;
3719: data <= 32'Hfffffffa;
3720: data <= 32'Hffffffff;
3721: data <= 32'H00000000;
3722: data <= 32'H00000008;
3723: data <= 32'H0000000f;
3724: data <= 32'H00000015;
3725: data <= 32'H00000010;
3726: data <= 32'H00000008;
3727: data <= 32'H00000003;
3728: data <= 32'H00000003;
3729: data <= 32'H00000005;
3730: data <= 32'H00000002;
3731: data <= 32'H00000000;
3732: data <= 32'H00000002;
3733: data <= 32'H00000002;
3734: data <= 32'H00000000;
3735: data <= 32'Hfffffffc;
3736: data <= 32'Hfffffffa;
3737: data <= 32'Hfffffff9;
3738: data <= 32'Hfffffffb;
3739: data <= 32'Hfffffff9;
3740: data <= 32'Hfffffff6;
3741: data <= 32'Hfffffff4;
3742: data <= 32'Hffffffef;
3743: data <= 32'Hffffffec;
3744: data <= 32'Hfffffff3;
3745: data <= 32'Hfffffff9;
3746: data <= 32'Hfffffff7;
3747: data <= 32'Hffffffed;
3748: data <= 32'Hffffffe7;
3749: data <= 32'Hffffffe5;
3750: data <= 32'Hffffffeb;
3751: data <= 32'Hffffffee;
3752: data <= 32'Hffffffef;
3753: data <= 32'Hfffffff2;
3754: data <= 32'Hfffffff5;
3755: data <= 32'Hfffffff4;
3756: data <= 32'Hfffffff1;
3757: data <= 32'Hffffffef;
3758: data <= 32'Hffffffe9;
3759: data <= 32'Hffffffec;
3760: data <= 32'Hffffffec;
3761: data <= 32'Hfffffff0;
3762: data <= 32'Hfffffff4;
3763: data <= 32'Hfffffff5;
3764: data <= 32'Hfffffffc;
3765: data <= 32'H00000004;
3766: data <= 32'H00000008;
3767: data <= 32'H00000009;
3768: data <= 32'H00000007;
3769: data <= 32'H00000002;
3770: data <= 32'H00000000;
3771: data <= 32'Hffffffff;
3772: data <= 32'Hffffffff;
3773: data <= 32'Hfffffffd;
3774: data <= 32'Hfffffffd;
3775: data <= 32'Hfffffffa;
3776: data <= 32'Hfffffffa;
3777: data <= 32'Hfffffff8;
3778: data <= 32'Hfffffff7;
3779: data <= 32'Hfffffff5;
3780: data <= 32'Hfffffff5;
3781: data <= 32'Hfffffff5;
3782: data <= 32'Hfffffff3;
3783: data <= 32'Hfffffff2;
3784: data <= 32'Hfffffff2;
3785: data <= 32'Hfffffff4;
3786: data <= 32'Hfffffff9;
3787: data <= 32'Hfffffff8;
3788: data <= 32'Hfffffff9;
3789: data <= 32'Hfffffff8;
3790: data <= 32'Hfffffff8;
3791: data <= 32'Hfffffff5;
3792: data <= 32'Hfffffff6;
3793: data <= 32'Hfffffff3;
3794: data <= 32'Hfffffff3;
3795: data <= 32'Hfffffff5;
3796: data <= 32'Hfffffff5;
3797: data <= 32'Hfffffff4;
3798: data <= 32'Hfffffff7;
3799: data <= 32'Hfffffff7;
3800: data <= 32'Hfffffff6;
3801: data <= 32'Hfffffff4;
3802: data <= 32'Hfffffff1;
3803: data <= 32'Hfffffff2;
3804: data <= 32'Hfffffff0;
3805: data <= 32'Hffffffef;
3806: data <= 32'Hffffffec;
3807: data <= 32'Hffffffee;
3808: data <= 32'Hffffffee;
3809: data <= 32'Hffffffec;
3810: data <= 32'Hffffffed;
3811: data <= 32'Hffffffea;
3812: data <= 32'Hffffffeb;
3813: data <= 32'Hffffffee;
3814: data <= 32'Hffffffed;
3815: data <= 32'Hfffffff1;
3816: data <= 32'Hffffffec;
3817: data <= 32'Hffffffed;
3818: data <= 32'Hffffffee;
3819: data <= 32'Hffffffed;
3820: data <= 32'Hfffffff1;
3821: data <= 32'Hfffffff9;
3822: data <= 32'Hfffffff7;
3823: data <= 32'Hfffffff8;
3824: data <= 32'Hfffffff6;
3825: data <= 32'Hfffffff9;
3826: data <= 32'H00000005;
3827: data <= 32'H00000009;
3828: data <= 32'H00000009;
3829: data <= 32'H0000000a;
3830: data <= 32'H00000006;
3831: data <= 32'Hffffffff;
3832: data <= 32'Hfffffffe;
3833: data <= 32'Hfffffff8;
3834: data <= 32'Hfffffff7;
3835: data <= 32'Hffffffff;
3836: data <= 32'H00000003;
3837: data <= 32'H00000000;
3838: data <= 32'Hfffffff5;
3839: data <= 32'Hffffffe9;
3840: data <= 32'Hffffffdf;
3841: data <= 32'Hfffffff4;
3842: data <= 32'Hfffffff1;
3843: data <= 32'Hfffffff3;
3844: data <= 32'Hfffffff4;
3845: data <= 32'Hfffffff1;
3846: data <= 32'Hfffffff0;
3847: data <= 32'Hfffffff3;
3848: data <= 32'Hfffffff7;
3849: data <= 32'Hfffffffa;
3850: data <= 32'Hfffffffc;
3851: data <= 32'H00000006;
3852: data <= 32'H0000000b;
3853: data <= 32'H00000006;
3854: data <= 32'H00000003;
3855: data <= 32'H00000002;
3856: data <= 32'Hffffffff;
3857: data <= 32'Hfffffffe;
3858: data <= 32'Hfffffffa;
3859: data <= 32'Hfffffff4;
3860: data <= 32'Hfffffff6;
3861: data <= 32'Hfffffff8;
3862: data <= 32'Hfffffff2;
3863: data <= 32'Hfffffff1;
3864: data <= 32'Hffffffef;
3865: data <= 32'Hffffffec;
3866: data <= 32'Hffffffec;
3867: data <= 32'Hffffffeb;
3868: data <= 32'Hffffffe6;
3869: data <= 32'Hffffffe4;
3870: data <= 32'Hffffffe4;
3871: data <= 32'Hffffffe6;
3872: data <= 32'Hfffffff2;
3873: data <= 32'Hfffffff9;
3874: data <= 32'Hfffffff7;
3875: data <= 32'Hffffffeb;
3876: data <= 32'Hffffffe4;
3877: data <= 32'Hffffffe4;
3878: data <= 32'Hffffffe8;
3879: data <= 32'Hffffffeb;
3880: data <= 32'Hffffffed;
3881: data <= 32'Hffffffed;
3882: data <= 32'Hffffffeb;
3883: data <= 32'Hffffffea;
3884: data <= 32'Hffffffe2;
3885: data <= 32'Hffffffdf;
3886: data <= 32'Hffffffda;
3887: data <= 32'Hffffffd7;
3888: data <= 32'Hffffffdc;
3889: data <= 32'Hffffffe5;
3890: data <= 32'Hffffffe9;
3891: data <= 32'Hffffffea;
3892: data <= 32'Hfffffff4;
3893: data <= 32'Hfffffffb;
3894: data <= 32'H00000003;
3895: data <= 32'H00000006;
3896: data <= 32'H00000002;
3897: data <= 32'H00000000;
3898: data <= 32'H00000000;
3899: data <= 32'Hfffffffc;
3900: data <= 32'Hfffffffa;
3901: data <= 32'Hfffffff8;
3902: data <= 32'Hfffffff7;
3903: data <= 32'Hfffffff7;
3904: data <= 32'Hfffffff5;
3905: data <= 32'Hfffffff3;
3906: data <= 32'Hfffffff0;
3907: data <= 32'Hfffffff2;
3908: data <= 32'Hffffffed;
3909: data <= 32'Hffffffee;
3910: data <= 32'Hffffffee;
3911: data <= 32'Hffffffea;
3912: data <= 32'Hffffffed;
3913: data <= 32'Hfffffff1;
3914: data <= 32'Hfffffff1;
3915: data <= 32'Hfffffff2;
3916: data <= 32'Hfffffff5;
3917: data <= 32'Hfffffff5;
3918: data <= 32'Hfffffff6;
3919: data <= 32'Hfffffff5;
3920: data <= 32'Hfffffff5;
3921: data <= 32'Hfffffff8;
3922: data <= 32'Hfffffff9;
3923: data <= 32'Hfffffffc;
3924: data <= 32'Hfffffffd;
3925: data <= 32'Hfffffffe;
3926: data <= 32'Hffffffff;
3927: data <= 32'Hfffffffb;
3928: data <= 32'Hfffffff8;
3929: data <= 32'Hfffffff3;
3930: data <= 32'Hfffffff0;
3931: data <= 32'Hfffffff1;
3932: data <= 32'Hffffffee;
3933: data <= 32'Hffffffea;
3934: data <= 32'Hffffffea;
3935: data <= 32'Hffffffe9;
3936: data <= 32'Hffffffe8;
3937: data <= 32'Hffffffe6;
3938: data <= 32'Hffffffe2;
3939: data <= 32'Hffffffe0;
3940: data <= 32'Hffffffe2;
3941: data <= 32'Hffffffe0;
3942: data <= 32'Hffffffe6;
3943: data <= 32'Hffffffe7;
3944: data <= 32'Hffffffe5;
3945: data <= 32'Hffffffe5;
3946: data <= 32'Hffffffe6;
3947: data <= 32'Hffffffe9;
3948: data <= 32'Hffffffec;
3949: data <= 32'Hfffffff3;
3950: data <= 32'Hfffffff7;
3951: data <= 32'Hfffffff3;
3952: data <= 32'Hffffffed;
3953: data <= 32'Hfffffff2;
3954: data <= 32'Hfffffff6;
3955: data <= 32'Hfffffffc;
3956: data <= 32'H00000000;
3957: data <= 32'Hfffffffd;
3958: data <= 32'H00000000;
3959: data <= 32'Hfffffffc;
3960: data <= 32'Hfffffff2;
3961: data <= 32'Hfffffff1;
3962: data <= 32'Hfffffff1;
3963: data <= 32'Hfffffff5;
3964: data <= 32'Hfffffffe;
3965: data <= 32'Hfffffffb;
3966: data <= 32'Hffffffeb;
3967: data <= 32'Hffffffe0;
3968: data <= 32'Hffffffd8;
3969: data <= 32'Hfffffff6;
3970: data <= 32'Hfffffff7;
3971: data <= 32'Hfffffff4;
3972: data <= 32'Hfffffff3;
3973: data <= 32'Hfffffff6;
3974: data <= 32'Hfffffff4;
3975: data <= 32'Hfffffff7;
3976: data <= 32'Hfffffff9;
3977: data <= 32'Hfffffffa;
3978: data <= 32'Hfffffffb;
3979: data <= 32'H00000001;
3980: data <= 32'H00000004;
3981: data <= 32'H00000001;
3982: data <= 32'H00000000;
3983: data <= 32'H00000003;
3984: data <= 32'H00000002;
3985: data <= 32'H00000002;
3986: data <= 32'Hfffffffc;
3987: data <= 32'Hfffffff5;
3988: data <= 32'Hfffffff6;
3989: data <= 32'Hfffffff5;
3990: data <= 32'Hfffffff5;
3991: data <= 32'Hfffffff1;
3992: data <= 32'Hffffffeb;
3993: data <= 32'Hffffffec;
3994: data <= 32'Hffffffea;
3995: data <= 32'Hffffffeb;
3996: data <= 32'Hffffffe8;
3997: data <= 32'Hffffffe1;
3998: data <= 32'Hffffffdf;
3999: data <= 32'Hffffffe1;
4000: data <= 32'Hfffffff2;
4001: data <= 32'Hfffffff9;
4002: data <= 32'Hfffffff7;
4003: data <= 32'Hfffffff2;
4004: data <= 32'Hffffffe9;
4005: data <= 32'Hffffffec;
4006: data <= 32'Hfffffff1;
4007: data <= 32'Hfffffff0;
4008: data <= 32'Hfffffff1;
4009: data <= 32'Hffffffef;
4010: data <= 32'Hffffffea;
4011: data <= 32'Hffffffe7;
4012: data <= 32'Hffffffe3;
4013: data <= 32'Hffffffd8;
4014: data <= 32'Hffffffd1;
4015: data <= 32'Hffffffce;
4016: data <= 32'Hffffffd2;
4017: data <= 32'Hffffffe0;
4018: data <= 32'Hffffffe4;
4019: data <= 32'Hffffffe9;
4020: data <= 32'Hfffffff1;
4021: data <= 32'Hfffffffa;
4022: data <= 32'H00000002;
4023: data <= 32'H00000004;
4024: data <= 32'H00000004;
4025: data <= 32'H00000002;
4026: data <= 32'H00000001;
4027: data <= 32'H00000001;
4028: data <= 32'Hfffffffc;
4029: data <= 32'Hfffffffb;
4030: data <= 32'Hfffffffc;
4031: data <= 32'Hfffffffa;
4032: data <= 32'Hfffffff9;
4033: data <= 32'Hfffffff7;
4034: data <= 32'Hfffffff8;
4035: data <= 32'Hfffffff7;
4036: data <= 32'Hfffffff4;
4037: data <= 32'Hfffffff5;
4038: data <= 32'Hfffffff0;
4039: data <= 32'Hfffffff3;
4040: data <= 32'Hfffffff4;
4041: data <= 32'Hfffffff2;
4042: data <= 32'Hfffffff4;
4043: data <= 32'Hfffffff3;
4044: data <= 32'Hfffffff4;
4045: data <= 32'Hfffffff6;
4046: data <= 32'Hfffffff5;
4047: data <= 32'Hfffffff6;
4048: data <= 32'Hfffffff8;
4049: data <= 32'Hfffffffd;
4050: data <= 32'Hfffffffc;
4051: data <= 32'H00000002;
4052: data <= 32'H00000001;
4053: data <= 32'H00000001;
4054: data <= 32'H00000002;
4055: data <= 32'Hfffffffb;
4056: data <= 32'Hfffffffa;
4057: data <= 32'Hfffffff8;
4058: data <= 32'Hfffffff0;
4059: data <= 32'Hffffffef;
4060: data <= 32'Hffffffed;
4061: data <= 32'Hffffffe9;
4062: data <= 32'Hffffffe8;
4063: data <= 32'Hffffffe7;
4064: data <= 32'Hffffffe5;
4065: data <= 32'Hffffffe2;
4066: data <= 32'Hffffffe4;
4067: data <= 32'Hffffffde;
4068: data <= 32'Hffffffde;
4069: data <= 32'Hffffffe1;
4070: data <= 32'Hffffffe2;
4071: data <= 32'Hffffffe2;
4072: data <= 32'Hffffffe1;
4073: data <= 32'Hffffffe1;
4074: data <= 32'Hffffffe5;
4075: data <= 32'Hffffffe8;
4076: data <= 32'Hffffffec;
4077: data <= 32'Hfffffff2;
4078: data <= 32'Hfffffff3;
4079: data <= 32'Hfffffff2;
4080: data <= 32'Hffffffed;
4081: data <= 32'Hffffffea;
4082: data <= 32'Hfffffff0;
4083: data <= 32'Hfffffff6;
4084: data <= 32'Hfffffff8;
4085: data <= 32'Hfffffff8;
4086: data <= 32'Hfffffffc;
4087: data <= 32'Hfffffffa;
4088: data <= 32'Hfffffff6;
4089: data <= 32'Hfffffff3;
4090: data <= 32'Hfffffff2;
4091: data <= 32'Hfffffff8;
4092: data <= 32'Hfffffff9;
4093: data <= 32'Hfffffff6;
4094: data <= 32'Hffffffea;
4095: data <= 32'Hffffffe1;
4096: data <= 32'Hffffffde;
4097: data <= 32'H00000003;
4098: data <= 32'H00000005;
4099: data <= 32'H00000002;
4100: data <= 32'H00000000;
4101: data <= 32'Hfffffffe;
4102: data <= 32'Hfffffffd;
4103: data <= 32'H00000000;
4104: data <= 32'H00000003;
4105: data <= 32'H00000001;
4106: data <= 32'H00000004;
4107: data <= 32'H00000007;
4108: data <= 32'H00000005;
4109: data <= 32'H00000002;
4110: data <= 32'H00000004;
4111: data <= 32'H00000009;
4112: data <= 32'H00000011;
4113: data <= 32'H0000000e;
4114: data <= 32'H0000000d;
4115: data <= 32'H00000005;
4116: data <= 32'H00000002;
4117: data <= 32'H00000005;
4118: data <= 32'H00000003;
4119: data <= 32'Hfffffffe;
4120: data <= 32'Hfffffff8;
4121: data <= 32'Hfffffff1;
4122: data <= 32'Hfffffff1;
4123: data <= 32'Hfffffff3;
4124: data <= 32'Hfffffff0;
4125: data <= 32'Hffffffe6;
4126: data <= 32'Hffffffde;
4127: data <= 32'Hffffffe4;
4128: data <= 32'Hfffffff1;
4129: data <= 32'Hfffffffb;
4130: data <= 32'Hfffffff8;
4131: data <= 32'Hfffffff1;
4132: data <= 32'Hffffffec;
4133: data <= 32'Hffffffeb;
4134: data <= 32'Hffffffeb;
4135: data <= 32'Hfffffff2;
4136: data <= 32'Hffffffed;
4137: data <= 32'Hffffffec;
4138: data <= 32'Hffffffea;
4139: data <= 32'Hffffffe7;
4140: data <= 32'Hffffffe6;
4141: data <= 32'Hffffffda;
4142: data <= 32'Hffffffd3;
4143: data <= 32'Hffffffd1;
4144: data <= 32'Hffffffd6;
4145: data <= 32'Hffffffe0;
4146: data <= 32'Hffffffe9;
4147: data <= 32'Hffffffea;
4148: data <= 32'Hfffffff6;
4149: data <= 32'Hffffffff;
4150: data <= 32'Hffffffff;
4151: data <= 32'H00000003;
4152: data <= 32'H00000004;
4153: data <= 32'H00000002;
4154: data <= 32'H00000002;
4155: data <= 32'H00000002;
4156: data <= 32'H00000000;
4157: data <= 32'Hffffffff;
4158: data <= 32'H00000000;
4159: data <= 32'H00000000;
4160: data <= 32'H00000001;
4161: data <= 32'Hfffffffe;
4162: data <= 32'H00000000;
4163: data <= 32'H00000001;
4164: data <= 32'Hfffffffa;
4165: data <= 32'Hfffffffa;
4166: data <= 32'Hfffffffb;
4167: data <= 32'Hfffffffc;
4168: data <= 32'Hfffffffc;
4169: data <= 32'Hfffffffc;
4170: data <= 32'Hfffffffa;
4171: data <= 32'Hfffffffa;
4172: data <= 32'Hfffffff8;
4173: data <= 32'Hfffffffa;
4174: data <= 32'Hfffffffb;
4175: data <= 32'Hfffffff9;
4176: data <= 32'Hfffffffc;
4177: data <= 32'Hffffffff;
4178: data <= 32'Hfffffffc;
4179: data <= 32'H00000000;
4180: data <= 32'H00000002;
4181: data <= 32'H00000002;
4182: data <= 32'Hfffffffe;
4183: data <= 32'Hfffffffe;
4184: data <= 32'Hfffffffa;
4185: data <= 32'Hfffffff7;
4186: data <= 32'Hfffffff2;
4187: data <= 32'Hffffffee;
4188: data <= 32'Hffffffe8;
4189: data <= 32'Hffffffe5;
4190: data <= 32'Hffffffe6;
4191: data <= 32'Hffffffe6;
4192: data <= 32'Hffffffe2;
4193: data <= 32'Hffffffe4;
4194: data <= 32'Hffffffe3;
4195: data <= 32'Hffffffe2;
4196: data <= 32'Hffffffe1;
4197: data <= 32'Hffffffe2;
4198: data <= 32'Hffffffe4;
4199: data <= 32'Hffffffe4;
4200: data <= 32'Hffffffe5;
4201: data <= 32'Hffffffe5;
4202: data <= 32'Hffffffea;
4203: data <= 32'Hffffffeb;
4204: data <= 32'Hffffffef;
4205: data <= 32'Hfffffff4;
4206: data <= 32'Hfffffff5;
4207: data <= 32'Hfffffff2;
4208: data <= 32'Hffffffef;
4209: data <= 32'Hffffffec;
4210: data <= 32'Hfffffff0;
4211: data <= 32'Hfffffff5;
4212: data <= 32'Hfffffff8;
4213: data <= 32'Hfffffff9;
4214: data <= 32'Hfffffffc;
4215: data <= 32'Hffffffff;
4216: data <= 32'Hfffffffd;
4217: data <= 32'Hfffffffb;
4218: data <= 32'Hfffffffa;
4219: data <= 32'Hfffffffd;
4220: data <= 32'H00000000;
4221: data <= 32'Hfffffffe;
4222: data <= 32'Hfffffff2;
4223: data <= 32'Hffffffee;
4224: data <= 32'Hffffffef;
4225: data <= 32'H0000000f;
4226: data <= 32'H0000000f;
4227: data <= 32'H0000000f;
4228: data <= 32'H0000000a;
4229: data <= 32'H00000007;
4230: data <= 32'H00000005;
4231: data <= 32'H00000006;
4232: data <= 32'H00000008;
4233: data <= 32'H0000000a;
4234: data <= 32'H00000009;
4235: data <= 32'H00000008;
4236: data <= 32'H00000008;
4237: data <= 32'Hfffffffc;
4238: data <= 32'H00000000;
4239: data <= 32'H0000000b;
4240: data <= 32'H00000013;
4241: data <= 32'H00000016;
4242: data <= 32'H0000000f;
4243: data <= 32'H00000008;
4244: data <= 32'H00000008;
4245: data <= 32'H00000007;
4246: data <= 32'H0000000b;
4247: data <= 32'H0000000c;
4248: data <= 32'H00000003;
4249: data <= 32'Hfffffffd;
4250: data <= 32'Hfffffffb;
4251: data <= 32'Hfffffffa;
4252: data <= 32'Hfffffff6;
4253: data <= 32'Hffffffea;
4254: data <= 32'Hffffffe2;
4255: data <= 32'Hffffffe8;
4256: data <= 32'Hfffffff5;
4257: data <= 32'Hfffffffd;
4258: data <= 32'Hfffffffb;
4259: data <= 32'Hfffffff7;
4260: data <= 32'Hffffffea;
4261: data <= 32'Hffffffeb;
4262: data <= 32'Hffffffeb;
4263: data <= 32'Hffffffee;
4264: data <= 32'Hffffffeb;
4265: data <= 32'Hffffffec;
4266: data <= 32'Hffffffe7;
4267: data <= 32'Hffffffeb;
4268: data <= 32'Hffffffee;
4269: data <= 32'Hffffffe2;
4270: data <= 32'Hffffffda;
4271: data <= 32'Hffffffd3;
4272: data <= 32'Hffffffd7;
4273: data <= 32'Hffffffe2;
4274: data <= 32'Hffffffea;
4275: data <= 32'Hffffffed;
4276: data <= 32'Hfffffff4;
4277: data <= 32'Hfffffffa;
4278: data <= 32'Hffffffff;
4279: data <= 32'Hfffffffc;
4280: data <= 32'Hfffffffe;
4281: data <= 32'Hfffffffd;
4282: data <= 32'Hfffffffc;
4283: data <= 32'Hfffffffb;
4284: data <= 32'Hfffffffe;
4285: data <= 32'Hfffffffa;
4286: data <= 32'Hfffffffc;
4287: data <= 32'Hfffffffd;
4288: data <= 32'Hffffffff;
4289: data <= 32'Hfffffffc;
4290: data <= 32'Hfffffffc;
4291: data <= 32'Hfffffffb;
4292: data <= 32'Hfffffffb;
4293: data <= 32'Hfffffff9;
4294: data <= 32'Hfffffff9;
4295: data <= 32'Hffffffff;
4296: data <= 32'Hfffffffd;
4297: data <= 32'Hfffffffd;
4298: data <= 32'Hfffffffe;
4299: data <= 32'Hfffffffe;
4300: data <= 32'Hfffffffa;
4301: data <= 32'Hfffffffe;
4302: data <= 32'Hfffffffc;
4303: data <= 32'Hffffffff;
4304: data <= 32'Hffffffff;
4305: data <= 32'Hffffffff;
4306: data <= 32'H00000001;
4307: data <= 32'H00000004;
4308: data <= 32'H00000002;
4309: data <= 32'H00000001;
4310: data <= 32'H00000000;
4311: data <= 32'Hffffffff;
4312: data <= 32'Hfffffffb;
4313: data <= 32'Hfffffff8;
4314: data <= 32'Hffffffef;
4315: data <= 32'Hffffffec;
4316: data <= 32'Hffffffe8;
4317: data <= 32'Hffffffe8;
4318: data <= 32'Hffffffe4;
4319: data <= 32'Hffffffe9;
4320: data <= 32'Hffffffe7;
4321: data <= 32'Hffffffe5;
4322: data <= 32'Hffffffea;
4323: data <= 32'Hffffffe7;
4324: data <= 32'Hffffffe6;
4325: data <= 32'Hffffffe6;
4326: data <= 32'Hffffffe9;
4327: data <= 32'Hffffffe8;
4328: data <= 32'Hffffffe6;
4329: data <= 32'Hffffffe9;
4330: data <= 32'Hffffffea;
4331: data <= 32'Hffffffea;
4332: data <= 32'Hffffffef;
4333: data <= 32'Hfffffff3;
4334: data <= 32'Hfffffff7;
4335: data <= 32'Hfffffff0;
4336: data <= 32'Hffffffee;
4337: data <= 32'Hffffffee;
4338: data <= 32'Hffffffef;
4339: data <= 32'Hfffffff5;
4340: data <= 32'Hfffffff9;
4341: data <= 32'Hfffffffa;
4342: data <= 32'H00000001;
4343: data <= 32'H00000002;
4344: data <= 32'H00000004;
4345: data <= 32'H00000008;
4346: data <= 32'H00000004;
4347: data <= 32'H00000008;
4348: data <= 32'H0000000d;
4349: data <= 32'H0000000a;
4350: data <= 32'H00000004;
4351: data <= 32'H00000002;
4352: data <= 32'Hfffffffd;
4353: data <= 32'H00000019;
4354: data <= 32'H0000001a;
4355: data <= 32'H00000017;
4356: data <= 32'H00000016;
4357: data <= 32'H00000012;
4358: data <= 32'H0000000f;
4359: data <= 32'H00000010;
4360: data <= 32'H00000011;
4361: data <= 32'H0000000f;
4362: data <= 32'H00000013;
4363: data <= 32'H00000012;
4364: data <= 32'H0000000f;
4365: data <= 32'H00000007;
4366: data <= 32'H00000000;
4367: data <= 32'H00000002;
4368: data <= 32'H00000013;
4369: data <= 32'H0000000f;
4370: data <= 32'H00000010;
4371: data <= 32'H0000000a;
4372: data <= 32'H00000003;
4373: data <= 32'H0000000a;
4374: data <= 32'H0000000e;
4375: data <= 32'H0000000e;
4376: data <= 32'H0000000b;
4377: data <= 32'H00000002;
4378: data <= 32'H00000002;
4379: data <= 32'Hffffffff;
4380: data <= 32'Hfffffffb;
4381: data <= 32'Hfffffff4;
4382: data <= 32'Hffffffec;
4383: data <= 32'Hffffffee;
4384: data <= 32'Hfffffffa;
4385: data <= 32'H00000005;
4386: data <= 32'H00000000;
4387: data <= 32'Hfffffff9;
4388: data <= 32'Hfffffff1;
4389: data <= 32'Hffffffee;
4390: data <= 32'Hffffffee;
4391: data <= 32'Hfffffff2;
4392: data <= 32'Hfffffff0;
4393: data <= 32'Hfffffff1;
4394: data <= 32'Hfffffff0;
4395: data <= 32'Hfffffff2;
4396: data <= 32'Hfffffff6;
4397: data <= 32'Hfffffff2;
4398: data <= 32'Hffffffe8;
4399: data <= 32'Hffffffe2;
4400: data <= 32'Hffffffe2;
4401: data <= 32'Hffffffea;
4402: data <= 32'Hfffffff5;
4403: data <= 32'Hfffffff6;
4404: data <= 32'Hfffffff8;
4405: data <= 32'Hffffffff;
4406: data <= 32'Hfffffffe;
4407: data <= 32'Hfffffffe;
4408: data <= 32'Hffffffff;
4409: data <= 32'Hfffffffd;
4410: data <= 32'Hfffffffd;
4411: data <= 32'Hfffffffe;
4412: data <= 32'Hffffffff;
4413: data <= 32'Hfffffffb;
4414: data <= 32'Hfffffffc;
4415: data <= 32'Hfffffffc;
4416: data <= 32'Hfffffff9;
4417: data <= 32'Hfffffffc;
4418: data <= 32'Hfffffff8;
4419: data <= 32'Hfffffff8;
4420: data <= 32'Hfffffffa;
4421: data <= 32'Hfffffff9;
4422: data <= 32'Hfffffffa;
4423: data <= 32'Hfffffffb;
4424: data <= 32'Hfffffffc;
4425: data <= 32'Hffffffff;
4426: data <= 32'Hffffffff;
4427: data <= 32'H00000001;
4428: data <= 32'Hffffffff;
4429: data <= 32'H00000000;
4430: data <= 32'H00000001;
4431: data <= 32'H00000003;
4432: data <= 32'H00000005;
4433: data <= 32'H00000005;
4434: data <= 32'H00000007;
4435: data <= 32'H0000000b;
4436: data <= 32'H00000007;
4437: data <= 32'H00000005;
4438: data <= 32'H00000004;
4439: data <= 32'H00000004;
4440: data <= 32'Hfffffffe;
4441: data <= 32'Hfffffffc;
4442: data <= 32'Hfffffff5;
4443: data <= 32'Hfffffff1;
4444: data <= 32'Hfffffff0;
4445: data <= 32'Hffffffee;
4446: data <= 32'Hffffffeb;
4447: data <= 32'Hffffffef;
4448: data <= 32'Hffffffef;
4449: data <= 32'Hffffffee;
4450: data <= 32'Hffffffef;
4451: data <= 32'Hffffffef;
4452: data <= 32'Hffffffef;
4453: data <= 32'Hffffffee;
4454: data <= 32'Hfffffff0;
4455: data <= 32'Hffffffee;
4456: data <= 32'Hfffffff3;
4457: data <= 32'Hfffffff2;
4458: data <= 32'Hfffffff4;
4459: data <= 32'Hfffffff1;
4460: data <= 32'Hfffffff8;
4461: data <= 32'Hfffffffb;
4462: data <= 32'Hfffffff8;
4463: data <= 32'Hfffffff8;
4464: data <= 32'Hfffffff5;
4465: data <= 32'Hfffffff1;
4466: data <= 32'Hfffffff4;
4467: data <= 32'Hfffffff8;
4468: data <= 32'Hfffffffa;
4469: data <= 32'H00000002;
4470: data <= 32'H00000001;
4471: data <= 32'H00000008;
4472: data <= 32'H0000000a;
4473: data <= 32'H0000000c;
4474: data <= 32'H00000010;
4475: data <= 32'H00000014;
4476: data <= 32'H00000017;
4477: data <= 32'H00000015;
4478: data <= 32'H00000012;
4479: data <= 32'H0000000e;
4480: data <= 32'H0000000d;
4481: data <= 32'H00000017;
4482: data <= 32'H00000016;
4483: data <= 32'H00000016;
4484: data <= 32'H00000015;
4485: data <= 32'H00000011;
4486: data <= 32'H00000011;
4487: data <= 32'H00000010;
4488: data <= 32'H00000010;
4489: data <= 32'H0000000f;
4490: data <= 32'H00000012;
4491: data <= 32'H0000000f;
4492: data <= 32'H00000012;
4493: data <= 32'H00000007;
4494: data <= 32'H00000002;
4495: data <= 32'Hffffffff;
4496: data <= 32'H00000004;
4497: data <= 32'H0000000a;
4498: data <= 32'H00000009;
4499: data <= 32'H00000006;
4500: data <= 32'H00000004;
4501: data <= 32'H00000007;
4502: data <= 32'H0000000b;
4503: data <= 32'H0000000c;
4504: data <= 32'H00000003;
4505: data <= 32'Hfffffffc;
4506: data <= 32'Hfffffffd;
4507: data <= 32'Hfffffffe;
4508: data <= 32'Hfffffff9;
4509: data <= 32'Hfffffff7;
4510: data <= 32'Hffffffee;
4511: data <= 32'Hffffffef;
4512: data <= 32'Hfffffff8;
4513: data <= 32'H00000004;
4514: data <= 32'H00000001;
4515: data <= 32'Hfffffffb;
4516: data <= 32'Hfffffff1;
4517: data <= 32'Hfffffff1;
4518: data <= 32'Hffffffee;
4519: data <= 32'Hffffffed;
4520: data <= 32'Hffffffef;
4521: data <= 32'Hffffffef;
4522: data <= 32'Hffffffec;
4523: data <= 32'Hffffffee;
4524: data <= 32'Hfffffff4;
4525: data <= 32'Hfffffff1;
4526: data <= 32'Hffffffec;
4527: data <= 32'Hffffffe4;
4528: data <= 32'Hffffffe4;
4529: data <= 32'Hffffffef;
4530: data <= 32'Hfffffff4;
4531: data <= 32'Hfffffffa;
4532: data <= 32'Hfffffff9;
4533: data <= 32'Hfffffffb;
4534: data <= 32'Hfffffffb;
4535: data <= 32'Hfffffff9;
4536: data <= 32'Hfffffffa;
4537: data <= 32'Hfffffffc;
4538: data <= 32'Hfffffffc;
4539: data <= 32'Hfffffffc;
4540: data <= 32'Hfffffffb;
4541: data <= 32'Hfffffff8;
4542: data <= 32'Hfffffff6;
4543: data <= 32'Hfffffff5;
4544: data <= 32'Hfffffff5;
4545: data <= 32'Hfffffff5;
4546: data <= 32'Hfffffff6;
4547: data <= 32'Hfffffff3;
4548: data <= 32'Hfffffff2;
4549: data <= 32'Hfffffff6;
4550: data <= 32'Hfffffff5;
4551: data <= 32'Hfffffff8;
4552: data <= 32'Hfffffff8;
4553: data <= 32'Hfffffffb;
4554: data <= 32'Hfffffffa;
4555: data <= 32'Hfffffffc;
4556: data <= 32'Hfffffffd;
4557: data <= 32'H00000002;
4558: data <= 32'H00000001;
4559: data <= 32'H00000005;
4560: data <= 32'H00000004;
4561: data <= 32'H00000008;
4562: data <= 32'H00000009;
4563: data <= 32'H0000000b;
4564: data <= 32'H00000007;
4565: data <= 32'H00000007;
4566: data <= 32'H00000005;
4567: data <= 32'H00000004;
4568: data <= 32'Hfffffffe;
4569: data <= 32'Hfffffff8;
4570: data <= 32'Hfffffff2;
4571: data <= 32'Hfffffff1;
4572: data <= 32'Hffffffee;
4573: data <= 32'Hffffffec;
4574: data <= 32'Hffffffee;
4575: data <= 32'Hffffffed;
4576: data <= 32'Hfffffff0;
4577: data <= 32'Hffffffed;
4578: data <= 32'Hfffffff0;
4579: data <= 32'Hfffffff3;
4580: data <= 32'Hfffffff1;
4581: data <= 32'Hfffffff0;
4582: data <= 32'Hffffffee;
4583: data <= 32'Hfffffff0;
4584: data <= 32'Hfffffff1;
4585: data <= 32'Hfffffff3;
4586: data <= 32'Hfffffff1;
4587: data <= 32'Hfffffff3;
4588: data <= 32'Hfffffff3;
4589: data <= 32'Hfffffff2;
4590: data <= 32'Hfffffff1;
4591: data <= 32'Hffffffeb;
4592: data <= 32'Hffffffeb;
4593: data <= 32'Hffffffec;
4594: data <= 32'Hffffffec;
4595: data <= 32'Hfffffff1;
4596: data <= 32'Hfffffff2;
4597: data <= 32'Hfffffff2;
4598: data <= 32'Hfffffff8;
4599: data <= 32'Hfffffffc;
4600: data <= 32'Hffffffff;
4601: data <= 32'H00000007;
4602: data <= 32'H0000000c;
4603: data <= 32'H00000010;
4604: data <= 32'H00000019;
4605: data <= 32'H00000013;
4606: data <= 32'H00000011;
4607: data <= 32'H00000010;
4608: data <= 32'H00000007;
4609: data <= 32'H00000011;
4610: data <= 32'H00000010;
4611: data <= 32'H00000010;
4612: data <= 32'H00000010;
4613: data <= 32'H0000000e;
4614: data <= 32'H0000000c;
4615: data <= 32'H0000000c;
4616: data <= 32'H0000000c;
4617: data <= 32'H0000000a;
4618: data <= 32'H0000000c;
4619: data <= 32'H0000000b;
4620: data <= 32'H00000009;
4621: data <= 32'H00000006;
4622: data <= 32'H00000001;
4623: data <= 32'Hfffffffc;
4624: data <= 32'H00000003;
4625: data <= 32'H00000002;
4626: data <= 32'H00000006;
4627: data <= 32'H00000009;
4628: data <= 32'H00000004;
4629: data <= 32'H00000007;
4630: data <= 32'H00000009;
4631: data <= 32'H00000009;
4632: data <= 32'H00000005;
4633: data <= 32'Hfffffffe;
4634: data <= 32'Hfffffffb;
4635: data <= 32'Hfffffffd;
4636: data <= 32'Hfffffffb;
4637: data <= 32'Hfffffff8;
4638: data <= 32'Hffffffef;
4639: data <= 32'Hfffffff2;
4640: data <= 32'Hfffffff8;
4641: data <= 32'Hfffffffe;
4642: data <= 32'H00000002;
4643: data <= 32'Hfffffffd;
4644: data <= 32'Hfffffff4;
4645: data <= 32'Hffffffef;
4646: data <= 32'Hfffffff1;
4647: data <= 32'Hffffffed;
4648: data <= 32'Hffffffe9;
4649: data <= 32'Hffffffe8;
4650: data <= 32'Hffffffe9;
4651: data <= 32'Hffffffe7;
4652: data <= 32'Hffffffeb;
4653: data <= 32'Hffffffef;
4654: data <= 32'Hffffffea;
4655: data <= 32'Hffffffe7;
4656: data <= 32'Hffffffe4;
4657: data <= 32'Hffffffec;
4658: data <= 32'Hfffffff7;
4659: data <= 32'Hfffffffa;
4660: data <= 32'Hfffffff9;
4661: data <= 32'Hfffffff9;
4662: data <= 32'Hfffffff9;
4663: data <= 32'Hfffffffc;
4664: data <= 32'Hfffffffc;
4665: data <= 32'Hffffffff;
4666: data <= 32'Hffffffff;
4667: data <= 32'Hfffffffc;
4668: data <= 32'Hfffffff8;
4669: data <= 32'Hfffffff6;
4670: data <= 32'Hfffffff4;
4671: data <= 32'Hfffffff4;
4672: data <= 32'Hfffffff1;
4673: data <= 32'Hfffffff2;
4674: data <= 32'Hfffffff4;
4675: data <= 32'Hffffffef;
4676: data <= 32'Hfffffff0;
4677: data <= 32'Hfffffff3;
4678: data <= 32'Hfffffff4;
4679: data <= 32'Hfffffff4;
4680: data <= 32'Hfffffff6;
4681: data <= 32'Hfffffff6;
4682: data <= 32'Hfffffffa;
4683: data <= 32'Hfffffffa;
4684: data <= 32'Hfffffffd;
4685: data <= 32'H00000001;
4686: data <= 32'H00000005;
4687: data <= 32'H00000006;
4688: data <= 32'H00000008;
4689: data <= 32'H00000008;
4690: data <= 32'H0000000b;
4691: data <= 32'H0000000b;
4692: data <= 32'H00000008;
4693: data <= 32'H00000008;
4694: data <= 32'H00000008;
4695: data <= 32'H00000002;
4696: data <= 32'Hfffffffa;
4697: data <= 32'Hfffffff3;
4698: data <= 32'Hffffffef;
4699: data <= 32'Hffffffeb;
4700: data <= 32'Hffffffe8;
4701: data <= 32'Hffffffe9;
4702: data <= 32'Hffffffeb;
4703: data <= 32'Hffffffed;
4704: data <= 32'Hfffffff0;
4705: data <= 32'Hffffffef;
4706: data <= 32'Hffffffef;
4707: data <= 32'Hfffffff3;
4708: data <= 32'Hfffffff1;
4709: data <= 32'Hffffffef;
4710: data <= 32'Hffffffef;
4711: data <= 32'Hffffffed;
4712: data <= 32'Hffffffed;
4713: data <= 32'Hffffffec;
4714: data <= 32'Hffffffed;
4715: data <= 32'Hffffffe8;
4716: data <= 32'Hffffffe7;
4717: data <= 32'Hffffffe9;
4718: data <= 32'Hffffffe1;
4719: data <= 32'Hffffffe7;
4720: data <= 32'Hffffffe4;
4721: data <= 32'Hffffffe4;
4722: data <= 32'Hffffffe8;
4723: data <= 32'Hffffffe6;
4724: data <= 32'Hffffffe1;
4725: data <= 32'Hffffffe6;
4726: data <= 32'Hffffffe9;
4727: data <= 32'Hffffffee;
4728: data <= 32'Hfffffff4;
4729: data <= 32'Hfffffff8;
4730: data <= 32'H00000001;
4731: data <= 32'H00000006;
4732: data <= 32'H0000000d;
4733: data <= 32'H0000000e;
4734: data <= 32'H00000007;
4735: data <= 32'H00000000;
4736: data <= 32'H00000001;
4737: data <= 32'H0000000f;
4738: data <= 32'H0000000b;
4739: data <= 32'H0000000c;
4740: data <= 32'H0000000d;
4741: data <= 32'H0000000b;
4742: data <= 32'H0000000b;
4743: data <= 32'H0000000c;
4744: data <= 32'H00000009;
4745: data <= 32'H0000000c;
4746: data <= 32'H0000000a;
4747: data <= 32'H0000000a;
4748: data <= 32'H00000009;
4749: data <= 32'H00000003;
4750: data <= 32'H00000000;
4751: data <= 32'Hffffffff;
4752: data <= 32'Hfffffff9;
4753: data <= 32'Hffffffff;
4754: data <= 32'H00000003;
4755: data <= 32'H0000000c;
4756: data <= 32'H00000009;
4757: data <= 32'H00000006;
4758: data <= 32'H00000007;
4759: data <= 32'H00000006;
4760: data <= 32'H00000006;
4761: data <= 32'H00000004;
4762: data <= 32'Hfffffffc;
4763: data <= 32'Hfffffffb;
4764: data <= 32'Hfffffffd;
4765: data <= 32'Hfffffff9;
4766: data <= 32'Hfffffff8;
4767: data <= 32'Hfffffff4;
4768: data <= 32'Hfffffff3;
4769: data <= 32'Hfffffffb;
4770: data <= 32'H00000001;
4771: data <= 32'Hfffffffd;
4772: data <= 32'Hfffffff7;
4773: data <= 32'Hfffffff1;
4774: data <= 32'Hffffffec;
4775: data <= 32'Hffffffea;
4776: data <= 32'Hffffffe6;
4777: data <= 32'Hffffffe6;
4778: data <= 32'Hffffffe3;
4779: data <= 32'Hffffffe0;
4780: data <= 32'Hffffffe6;
4781: data <= 32'Hffffffee;
4782: data <= 32'Hffffffeb;
4783: data <= 32'Hffffffe7;
4784: data <= 32'Hffffffe2;
4785: data <= 32'Hffffffe8;
4786: data <= 32'Hffffffef;
4787: data <= 32'Hfffffffa;
4788: data <= 32'Hfffffff8;
4789: data <= 32'Hfffffff5;
4790: data <= 32'Hfffffff8;
4791: data <= 32'Hfffffffa;
4792: data <= 32'Hfffffffc;
4793: data <= 32'Hfffffffd;
4794: data <= 32'Hfffffffd;
4795: data <= 32'Hfffffff8;
4796: data <= 32'Hfffffff4;
4797: data <= 32'Hfffffff5;
4798: data <= 32'Hfffffff4;
4799: data <= 32'Hfffffff3;
4800: data <= 32'Hfffffff1;
4801: data <= 32'Hffffffee;
4802: data <= 32'Hffffffee;
4803: data <= 32'Hffffffec;
4804: data <= 32'Hffffffeb;
4805: data <= 32'Hffffffeb;
4806: data <= 32'Hffffffef;
4807: data <= 32'Hffffffef;
4808: data <= 32'Hfffffff1;
4809: data <= 32'Hfffffff5;
4810: data <= 32'Hfffffffa;
4811: data <= 32'Hfffffffa;
4812: data <= 32'H00000002;
4813: data <= 32'H00000002;
4814: data <= 32'H00000008;
4815: data <= 32'H00000007;
4816: data <= 32'H00000009;
4817: data <= 32'H0000000a;
4818: data <= 32'H0000000e;
4819: data <= 32'H0000000b;
4820: data <= 32'H00000008;
4821: data <= 32'H00000008;
4822: data <= 32'H00000008;
4823: data <= 32'H00000000;
4824: data <= 32'Hfffffff8;
4825: data <= 32'Hfffffff0;
4826: data <= 32'Hffffffeb;
4827: data <= 32'Hffffffeb;
4828: data <= 32'Hffffffe6;
4829: data <= 32'Hffffffe8;
4830: data <= 32'Hffffffeb;
4831: data <= 32'Hffffffe9;
4832: data <= 32'Hfffffff0;
4833: data <= 32'Hfffffff1;
4834: data <= 32'Hfffffff0;
4835: data <= 32'Hfffffff0;
4836: data <= 32'Hfffffff2;
4837: data <= 32'Hffffffed;
4838: data <= 32'Hffffffea;
4839: data <= 32'Hffffffeb;
4840: data <= 32'Hffffffe9;
4841: data <= 32'Hffffffe7;
4842: data <= 32'Hffffffe1;
4843: data <= 32'Hffffffdf;
4844: data <= 32'Hffffffdd;
4845: data <= 32'Hffffffde;
4846: data <= 32'Hffffffd9;
4847: data <= 32'Hffffffde;
4848: data <= 32'Hffffffde;
4849: data <= 32'Hffffffde;
4850: data <= 32'Hffffffdc;
4851: data <= 32'Hffffffdc;
4852: data <= 32'Hffffffd7;
4853: data <= 32'Hffffffda;
4854: data <= 32'Hffffffe1;
4855: data <= 32'Hffffffe5;
4856: data <= 32'Hffffffe9;
4857: data <= 32'Hffffffee;
4858: data <= 32'Hfffffff7;
4859: data <= 32'Hffffffff;
4860: data <= 32'H00000005;
4861: data <= 32'Hffffffff;
4862: data <= 32'Hfffffff9;
4863: data <= 32'Hfffffffa;
4864: data <= 32'Hfffffff8;
4865: data <= 32'H0000000b;
4866: data <= 32'H0000000d;
4867: data <= 32'H0000000c;
4868: data <= 32'H00000008;
4869: data <= 32'H00000012;
4870: data <= 32'H0000000d;
4871: data <= 32'H0000000c;
4872: data <= 32'H0000000e;
4873: data <= 32'H0000000f;
4874: data <= 32'H0000000d;
4875: data <= 32'H0000000f;
4876: data <= 32'H0000000e;
4877: data <= 32'H00000007;
4878: data <= 32'H00000003;
4879: data <= 32'Hfffffffc;
4880: data <= 32'Hfffffff6;
4881: data <= 32'Hfffffff8;
4882: data <= 32'Hfffffffd;
4883: data <= 32'H00000006;
4884: data <= 32'H0000000b;
4885: data <= 32'H00000009;
4886: data <= 32'H00000003;
4887: data <= 32'H00000004;
4888: data <= 32'H00000005;
4889: data <= 32'H00000003;
4890: data <= 32'Hfffffffe;
4891: data <= 32'Hfffffff5;
4892: data <= 32'Hfffffff6;
4893: data <= 32'Hfffffffa;
4894: data <= 32'Hfffffffe;
4895: data <= 32'Hfffffff5;
4896: data <= 32'Hfffffff1;
4897: data <= 32'Hfffffff1;
4898: data <= 32'Hfffffffb;
4899: data <= 32'Hffffffff;
4900: data <= 32'Hfffffff7;
4901: data <= 32'Hfffffff0;
4902: data <= 32'Hffffffea;
4903: data <= 32'Hffffffe4;
4904: data <= 32'Hffffffe4;
4905: data <= 32'Hffffffe5;
4906: data <= 32'Hffffffde;
4907: data <= 32'Hffffffdd;
4908: data <= 32'Hffffffe2;
4909: data <= 32'Hfffffff1;
4910: data <= 32'Hfffffff3;
4911: data <= 32'Hffffffef;
4912: data <= 32'Hffffffe7;
4913: data <= 32'Hffffffe6;
4914: data <= 32'Hffffffed;
4915: data <= 32'Hfffffff7;
4916: data <= 32'Hfffffff8;
4917: data <= 32'Hfffffff6;
4918: data <= 32'Hfffffff4;
4919: data <= 32'Hfffffff5;
4920: data <= 32'Hfffffff6;
4921: data <= 32'Hfffffff7;
4922: data <= 32'Hfffffff6;
4923: data <= 32'Hfffffff1;
4924: data <= 32'Hfffffff1;
4925: data <= 32'Hffffffef;
4926: data <= 32'Hfffffff0;
4927: data <= 32'Hffffffee;
4928: data <= 32'Hffffffee;
4929: data <= 32'Hffffffea;
4930: data <= 32'Hffffffe7;
4931: data <= 32'Hffffffe6;
4932: data <= 32'Hffffffe4;
4933: data <= 32'Hffffffe4;
4934: data <= 32'Hffffffe6;
4935: data <= 32'Hffffffe8;
4936: data <= 32'Hfffffff0;
4937: data <= 32'Hfffffff2;
4938: data <= 32'Hfffffffa;
4939: data <= 32'H00000000;
4940: data <= 32'H00000004;
4941: data <= 32'H00000007;
4942: data <= 32'H0000000b;
4943: data <= 32'H0000000a;
4944: data <= 32'H0000000c;
4945: data <= 32'H0000000c;
4946: data <= 32'H0000000e;
4947: data <= 32'H0000000a;
4948: data <= 32'H0000000a;
4949: data <= 32'H00000009;
4950: data <= 32'H00000009;
4951: data <= 32'H00000003;
4952: data <= 32'Hfffffff9;
4953: data <= 32'Hfffffff2;
4954: data <= 32'Hfffffff0;
4955: data <= 32'Hffffffeb;
4956: data <= 32'Hffffffe9;
4957: data <= 32'Hffffffe8;
4958: data <= 32'Hffffffea;
4959: data <= 32'Hffffffeb;
4960: data <= 32'Hffffffed;
4961: data <= 32'Hfffffff0;
4962: data <= 32'Hfffffff3;
4963: data <= 32'Hffffffef;
4964: data <= 32'Hfffffff1;
4965: data <= 32'Hffffffed;
4966: data <= 32'Hffffffeb;
4967: data <= 32'Hffffffea;
4968: data <= 32'Hffffffe8;
4969: data <= 32'Hffffffe2;
4970: data <= 32'Hffffffdd;
4971: data <= 32'Hffffffdc;
4972: data <= 32'Hffffffda;
4973: data <= 32'Hffffffdb;
4974: data <= 32'Hffffffd5;
4975: data <= 32'Hffffffd3;
4976: data <= 32'Hffffffd4;
4977: data <= 32'Hffffffd3;
4978: data <= 32'Hffffffd0;
4979: data <= 32'Hffffffd0;
4980: data <= 32'Hffffffd2;
4981: data <= 32'Hffffffd7;
4982: data <= 32'Hffffffdb;
4983: data <= 32'Hffffffe0;
4984: data <= 32'Hffffffe0;
4985: data <= 32'Hffffffe3;
4986: data <= 32'Hffffffec;
4987: data <= 32'Hfffffff4;
4988: data <= 32'Hfffffff4;
4989: data <= 32'Hfffffff1;
4990: data <= 32'Hfffffff0;
4991: data <= 32'Hfffffff1;
4992: data <= 32'Hfffffffa;
4993: data <= 32'H00000009;
4994: data <= 32'H00000006;
4995: data <= 32'H00000006;
4996: data <= 32'H00000008;
4997: data <= 32'H00000009;
4998: data <= 32'H00000008;
4999: data <= 32'H00000008;
5000: data <= 32'H00000009;
5001: data <= 32'H0000000a;
5002: data <= 32'H0000000b;
5003: data <= 32'H0000000b;
5004: data <= 32'H0000000b;
5005: data <= 32'H00000007;
5006: data <= 32'H00000001;
5007: data <= 32'Hfffffffb;
5008: data <= 32'Hfffffff1;
5009: data <= 32'Hfffffff0;
5010: data <= 32'Hfffffff1;
5011: data <= 32'Hfffffff9;
5012: data <= 32'H00000004;
5013: data <= 32'H00000007;
5014: data <= 32'H00000004;
5015: data <= 32'Hffffffff;
5016: data <= 32'H00000001;
5017: data <= 32'H00000000;
5018: data <= 32'Hfffffffa;
5019: data <= 32'Hfffffff3;
5020: data <= 32'Hfffffff0;
5021: data <= 32'Hfffffff1;
5022: data <= 32'Hfffffffb;
5023: data <= 32'Hfffffff4;
5024: data <= 32'Hffffffef;
5025: data <= 32'Hffffffe8;
5026: data <= 32'Hffffffee;
5027: data <= 32'Hfffffff4;
5028: data <= 32'Hfffffff3;
5029: data <= 32'Hffffffef;
5030: data <= 32'Hffffffe5;
5031: data <= 32'Hffffffe1;
5032: data <= 32'Hffffffdc;
5033: data <= 32'Hffffffdb;
5034: data <= 32'Hffffffdc;
5035: data <= 32'Hffffffd9;
5036: data <= 32'Hffffffdf;
5037: data <= 32'Hffffffeb;
5038: data <= 32'Hfffffff3;
5039: data <= 32'Hfffffffa;
5040: data <= 32'Hfffffff3;
5041: data <= 32'Hffffffe8;
5042: data <= 32'Hffffffe9;
5043: data <= 32'Hfffffff1;
5044: data <= 32'Hfffffff3;
5045: data <= 32'Hfffffff7;
5046: data <= 32'Hfffffff1;
5047: data <= 32'Hffffffec;
5048: data <= 32'Hffffffeb;
5049: data <= 32'Hffffffe9;
5050: data <= 32'Hffffffeb;
5051: data <= 32'Hffffffe7;
5052: data <= 32'Hffffffe5;
5053: data <= 32'Hffffffe5;
5054: data <= 32'Hffffffe5;
5055: data <= 32'Hffffffe4;
5056: data <= 32'Hffffffe6;
5057: data <= 32'Hffffffe4;
5058: data <= 32'Hffffffdf;
5059: data <= 32'Hffffffdc;
5060: data <= 32'Hffffffd8;
5061: data <= 32'Hffffffd8;
5062: data <= 32'Hffffffdb;
5063: data <= 32'Hffffffdd;
5064: data <= 32'Hffffffe1;
5065: data <= 32'Hffffffea;
5066: data <= 32'Hfffffff3;
5067: data <= 32'Hfffffff7;
5068: data <= 32'Hffffffff;
5069: data <= 32'Hfffffffe;
5070: data <= 32'Hffffffff;
5071: data <= 32'Hfffffffd;
5072: data <= 32'Hfffffffe;
5073: data <= 32'Hfffffffc;
5074: data <= 32'Hfffffffc;
5075: data <= 32'Hfffffffd;
5076: data <= 32'Hfffffffc;
5077: data <= 32'Hfffffffb;
5078: data <= 32'Hfffffffd;
5079: data <= 32'Hfffffff9;
5080: data <= 32'Hfffffff6;
5081: data <= 32'Hfffffff0;
5082: data <= 32'Hffffffec;
5083: data <= 32'Hffffffec;
5084: data <= 32'Hffffffe9;
5085: data <= 32'Hffffffe9;
5086: data <= 32'Hffffffe9;
5087: data <= 32'Hffffffe9;
5088: data <= 32'Hffffffe9;
5089: data <= 32'Hffffffe9;
5090: data <= 32'Hffffffed;
5091: data <= 32'Hffffffeb;
5092: data <= 32'Hffffffeb;
5093: data <= 32'Hffffffea;
5094: data <= 32'Hffffffe9;
5095: data <= 32'Hffffffe7;
5096: data <= 32'Hffffffe6;
5097: data <= 32'Hffffffe1;
5098: data <= 32'Hffffffdc;
5099: data <= 32'Hffffffdc;
5100: data <= 32'Hffffffd9;
5101: data <= 32'Hffffffd2;
5102: data <= 32'Hffffffcd;
5103: data <= 32'Hffffffc7;
5104: data <= 32'Hffffffc8;
5105: data <= 32'Hffffffca;
5106: data <= 32'Hffffffcd;
5107: data <= 32'Hffffffd1;
5108: data <= 32'Hffffffd8;
5109: data <= 32'Hffffffdc;
5110: data <= 32'Hffffffdb;
5111: data <= 32'Hffffffda;
5112: data <= 32'Hffffffdc;
5113: data <= 32'Hffffffdf;
5114: data <= 32'Hffffffe5;
5115: data <= 32'Hffffffe7;
5116: data <= 32'Hffffffe5;
5117: data <= 32'Hffffffe6;
5118: data <= 32'Hffffffea;
5119: data <= 32'Hfffffff4;
5120: data <= 32'Hfffffffe;
5121: data <= 32'H00000006;
5122: data <= 32'H00000004;
5123: data <= 32'H00000006;
5124: data <= 32'H00000008;
5125: data <= 32'H00000008;
5126: data <= 32'H00000006;
5127: data <= 32'H00000007;
5128: data <= 32'H00000007;
5129: data <= 32'H00000008;
5130: data <= 32'H00000009;
5131: data <= 32'H0000000a;
5132: data <= 32'H0000000b;
5133: data <= 32'H00000007;
5134: data <= 32'H00000005;
5135: data <= 32'H00000002;
5136: data <= 32'Hfffffff6;
5137: data <= 32'Hfffffff3;
5138: data <= 32'Hfffffff1;
5139: data <= 32'Hfffffff3;
5140: data <= 32'Hffffffff;
5141: data <= 32'H00000005;
5142: data <= 32'H00000009;
5143: data <= 32'H00000004;
5144: data <= 32'H00000002;
5145: data <= 32'H00000001;
5146: data <= 32'H00000002;
5147: data <= 32'Hfffffff8;
5148: data <= 32'Hfffffff1;
5149: data <= 32'Hfffffff4;
5150: data <= 32'Hfffffff7;
5151: data <= 32'Hfffffff9;
5152: data <= 32'Hfffffff7;
5153: data <= 32'Hfffffff1;
5154: data <= 32'Hffffffec;
5155: data <= 32'Hfffffff4;
5156: data <= 32'Hfffffff9;
5157: data <= 32'Hfffffff9;
5158: data <= 32'Hfffffff3;
5159: data <= 32'Hffffffe8;
5160: data <= 32'Hffffffe6;
5161: data <= 32'Hffffffe2;
5162: data <= 32'Hffffffe0;
5163: data <= 32'Hffffffe3;
5164: data <= 32'Hffffffe1;
5165: data <= 32'Hffffffe4;
5166: data <= 32'Hfffffff4;
5167: data <= 32'H00000000;
5168: data <= 32'H00000000;
5169: data <= 32'Hfffffff3;
5170: data <= 32'Hffffffeb;
5171: data <= 32'Hffffffec;
5172: data <= 32'Hfffffff4;
5173: data <= 32'Hfffffff8;
5174: data <= 32'Hfffffff0;
5175: data <= 32'Hffffffee;
5176: data <= 32'Hffffffe5;
5177: data <= 32'Hffffffe0;
5178: data <= 32'Hffffffde;
5179: data <= 32'Hffffffdf;
5180: data <= 32'Hffffffe2;
5181: data <= 32'Hffffffe0;
5182: data <= 32'Hffffffe1;
5183: data <= 32'Hffffffe2;
5184: data <= 32'Hffffffe1;
5185: data <= 32'Hffffffe2;
5186: data <= 32'Hffffffe1;
5187: data <= 32'Hffffffdc;
5188: data <= 32'Hffffffd9;
5189: data <= 32'Hffffffda;
5190: data <= 32'Hffffffd5;
5191: data <= 32'Hffffffd7;
5192: data <= 32'Hffffffdc;
5193: data <= 32'Hffffffe2;
5194: data <= 32'Hffffffeb;
5195: data <= 32'Hffffffef;
5196: data <= 32'Hfffffff1;
5197: data <= 32'Hfffffff5;
5198: data <= 32'Hfffffff2;
5199: data <= 32'Hfffffff2;
5200: data <= 32'Hffffffec;
5201: data <= 32'Hffffffe9;
5202: data <= 32'Hffffffed;
5203: data <= 32'Hffffffeb;
5204: data <= 32'Hffffffe9;
5205: data <= 32'Hffffffef;
5206: data <= 32'Hffffffef;
5207: data <= 32'Hfffffff0;
5208: data <= 32'Hfffffff1;
5209: data <= 32'Hffffffec;
5210: data <= 32'Hffffffee;
5211: data <= 32'Hfffffff0;
5212: data <= 32'Hfffffff0;
5213: data <= 32'Hffffffed;
5214: data <= 32'Hffffffee;
5215: data <= 32'Hffffffef;
5216: data <= 32'Hffffffec;
5217: data <= 32'Hffffffec;
5218: data <= 32'Hffffffec;
5219: data <= 32'Hffffffec;
5220: data <= 32'Hffffffeb;
5221: data <= 32'Hffffffec;
5222: data <= 32'Hffffffeb;
5223: data <= 32'Hffffffe9;
5224: data <= 32'Hffffffea;
5225: data <= 32'Hffffffe7;
5226: data <= 32'Hffffffe5;
5227: data <= 32'Hffffffe3;
5228: data <= 32'Hffffffd8;
5229: data <= 32'Hffffffcd;
5230: data <= 32'Hffffffcb;
5231: data <= 32'Hffffffcc;
5232: data <= 32'Hffffffd0;
5233: data <= 32'Hffffffd5;
5234: data <= 32'Hffffffdb;
5235: data <= 32'Hffffffe0;
5236: data <= 32'Hffffffe6;
5237: data <= 32'Hffffffe3;
5238: data <= 32'Hffffffe7;
5239: data <= 32'Hffffffe6;
5240: data <= 32'Hffffffe9;
5241: data <= 32'Hffffffe9;
5242: data <= 32'Hffffffe5;
5243: data <= 32'Hffffffea;
5244: data <= 32'Hffffffe9;
5245: data <= 32'Hffffffe8;
5246: data <= 32'Hfffffff1;
5247: data <= 32'Hfffffff9;
5248: data <= 32'Hfffffffd;
5249: data <= 32'H00000002;
5250: data <= 32'H00000003;
5251: data <= 32'H00000004;
5252: data <= 32'H00000007;
5253: data <= 32'H00000004;
5254: data <= 32'H00000004;
5255: data <= 32'H00000006;
5256: data <= 32'H00000005;
5257: data <= 32'H00000005;
5258: data <= 32'H00000008;
5259: data <= 32'H00000005;
5260: data <= 32'H00000004;
5261: data <= 32'H00000006;
5262: data <= 32'H00000005;
5263: data <= 32'H00000001;
5264: data <= 32'Hfffffffd;
5265: data <= 32'Hfffffff7;
5266: data <= 32'Hfffffff1;
5267: data <= 32'Hfffffff0;
5268: data <= 32'Hfffffff5;
5269: data <= 32'Hffffffff;
5270: data <= 32'H00000008;
5271: data <= 32'H00000004;
5272: data <= 32'H00000004;
5273: data <= 32'H00000003;
5274: data <= 32'H00000002;
5275: data <= 32'Hfffffffd;
5276: data <= 32'Hfffffff7;
5277: data <= 32'Hfffffff3;
5278: data <= 32'Hfffffff2;
5279: data <= 32'Hfffffff9;
5280: data <= 32'Hfffffffb;
5281: data <= 32'Hfffffff6;
5282: data <= 32'Hfffffff2;
5283: data <= 32'Hfffffff5;
5284: data <= 32'Hfffffffd;
5285: data <= 32'H00000002;
5286: data <= 32'Hfffffffd;
5287: data <= 32'Hfffffff7;
5288: data <= 32'Hfffffff1;
5289: data <= 32'Hffffffec;
5290: data <= 32'Hffffffed;
5291: data <= 32'Hffffffeb;
5292: data <= 32'Hffffffed;
5293: data <= 32'Hffffffec;
5294: data <= 32'Hfffffff1;
5295: data <= 32'Hfffffffe;
5296: data <= 32'H00000008;
5297: data <= 32'Hfffffffe;
5298: data <= 32'Hfffffff9;
5299: data <= 32'Hfffffff1;
5300: data <= 32'Hfffffff1;
5301: data <= 32'Hfffffff8;
5302: data <= 32'Hfffffff6;
5303: data <= 32'Hfffffff4;
5304: data <= 32'Hffffffe9;
5305: data <= 32'Hffffffe0;
5306: data <= 32'Hffffffd9;
5307: data <= 32'Hffffffde;
5308: data <= 32'Hffffffe2;
5309: data <= 32'Hffffffe4;
5310: data <= 32'Hffffffe5;
5311: data <= 32'Hffffffe6;
5312: data <= 32'Hffffffe6;
5313: data <= 32'Hffffffe7;
5314: data <= 32'Hffffffe4;
5315: data <= 32'Hffffffe1;
5316: data <= 32'Hffffffe0;
5317: data <= 32'Hffffffdb;
5318: data <= 32'Hffffffd8;
5319: data <= 32'Hffffffd8;
5320: data <= 32'Hffffffd8;
5321: data <= 32'Hffffffdb;
5322: data <= 32'Hffffffdf;
5323: data <= 32'Hffffffe4;
5324: data <= 32'Hffffffe5;
5325: data <= 32'Hffffffe9;
5326: data <= 32'Hffffffe9;
5327: data <= 32'Hffffffe6;
5328: data <= 32'Hffffffe1;
5329: data <= 32'Hffffffe1;
5330: data <= 32'Hffffffde;
5331: data <= 32'Hffffffdf;
5332: data <= 32'Hffffffdf;
5333: data <= 32'Hffffffe2;
5334: data <= 32'Hffffffe3;
5335: data <= 32'Hffffffe3;
5336: data <= 32'Hffffffe8;
5337: data <= 32'Hffffffe7;
5338: data <= 32'Hffffffea;
5339: data <= 32'Hffffffec;
5340: data <= 32'Hffffffef;
5341: data <= 32'Hffffffef;
5342: data <= 32'Hffffffed;
5343: data <= 32'Hfffffff0;
5344: data <= 32'Hfffffff0;
5345: data <= 32'Hffffffec;
5346: data <= 32'Hffffffef;
5347: data <= 32'Hffffffee;
5348: data <= 32'Hffffffed;
5349: data <= 32'Hffffffee;
5350: data <= 32'Hffffffec;
5351: data <= 32'Hffffffea;
5352: data <= 32'Hffffffec;
5353: data <= 32'Hffffffed;
5354: data <= 32'Hffffffe9;
5355: data <= 32'Hffffffe0;
5356: data <= 32'Hffffffdb;
5357: data <= 32'Hffffffd2;
5358: data <= 32'Hffffffd1;
5359: data <= 32'Hffffffda;
5360: data <= 32'Hffffffdd;
5361: data <= 32'Hffffffdf;
5362: data <= 32'Hffffffe7;
5363: data <= 32'Hffffffe7;
5364: data <= 32'Hffffffed;
5365: data <= 32'Hfffffff0;
5366: data <= 32'Hfffffff0;
5367: data <= 32'Hfffffff0;
5368: data <= 32'Hfffffff2;
5369: data <= 32'Hffffffef;
5370: data <= 32'Hfffffff2;
5371: data <= 32'Hfffffff1;
5372: data <= 32'Hffffffee;
5373: data <= 32'Hffffffef;
5374: data <= 32'Hfffffff1;
5375: data <= 32'Hfffffff8;
5376: data <= 32'Hffffffff;
5377: data <= 32'H00000006;
5378: data <= 32'H00000004;
5379: data <= 32'H00000003;
5380: data <= 32'H00000006;
5381: data <= 32'H00000004;
5382: data <= 32'H00000006;
5383: data <= 32'H00000007;
5384: data <= 32'H00000007;
5385: data <= 32'H00000008;
5386: data <= 32'H00000004;
5387: data <= 32'H00000004;
5388: data <= 32'H00000007;
5389: data <= 32'H00000006;
5390: data <= 32'H00000007;
5391: data <= 32'H00000006;
5392: data <= 32'H00000003;
5393: data <= 32'H00000000;
5394: data <= 32'Hfffffff7;
5395: data <= 32'Hfffffff2;
5396: data <= 32'Hfffffff4;
5397: data <= 32'Hfffffff7;
5398: data <= 32'H00000000;
5399: data <= 32'H00000006;
5400: data <= 32'H00000005;
5401: data <= 32'H00000007;
5402: data <= 32'H00000004;
5403: data <= 32'H00000001;
5404: data <= 32'Hfffffffc;
5405: data <= 32'Hfffffff7;
5406: data <= 32'Hfffffff3;
5407: data <= 32'Hfffffff5;
5408: data <= 32'Hfffffff7;
5409: data <= 32'Hfffffffa;
5410: data <= 32'Hfffffff6;
5411: data <= 32'Hfffffff9;
5412: data <= 32'Hfffffffc;
5413: data <= 32'H00000003;
5414: data <= 32'H00000008;
5415: data <= 32'H00000004;
5416: data <= 32'Hfffffffe;
5417: data <= 32'Hfffffff9;
5418: data <= 32'Hfffffff6;
5419: data <= 32'Hfffffff7;
5420: data <= 32'Hfffffffa;
5421: data <= 32'Hfffffff4;
5422: data <= 32'Hfffffff6;
5423: data <= 32'Hfffffffa;
5424: data <= 32'H00000007;
5425: data <= 32'H0000000d;
5426: data <= 32'H00000007;
5427: data <= 32'Hfffffffd;
5428: data <= 32'Hfffffff2;
5429: data <= 32'Hfffffff7;
5430: data <= 32'Hfffffffa;
5431: data <= 32'Hfffffff9;
5432: data <= 32'Hffffffed;
5433: data <= 32'Hffffffe4;
5434: data <= 32'Hffffffde;
5435: data <= 32'Hffffffdb;
5436: data <= 32'Hffffffe2;
5437: data <= 32'Hffffffe6;
5438: data <= 32'Hffffffeb;
5439: data <= 32'Hffffffec;
5440: data <= 32'Hffffffee;
5441: data <= 32'Hffffffee;
5442: data <= 32'Hffffffeb;
5443: data <= 32'Hffffffe8;
5444: data <= 32'Hffffffe6;
5445: data <= 32'Hffffffdf;
5446: data <= 32'Hffffffda;
5447: data <= 32'Hffffffdb;
5448: data <= 32'Hffffffd7;
5449: data <= 32'Hffffffd5;
5450: data <= 32'Hffffffd5;
5451: data <= 32'Hffffffdb;
5452: data <= 32'Hffffffe0;
5453: data <= 32'Hffffffe5;
5454: data <= 32'Hffffffdf;
5455: data <= 32'Hffffffdf;
5456: data <= 32'Hffffffdd;
5457: data <= 32'Hffffffdc;
5458: data <= 32'Hffffffdf;
5459: data <= 32'Hffffffe1;
5460: data <= 32'Hffffffde;
5461: data <= 32'Hffffffe1;
5462: data <= 32'Hffffffde;
5463: data <= 32'Hffffffe1;
5464: data <= 32'Hffffffe4;
5465: data <= 32'Hffffffe5;
5466: data <= 32'Hffffffe9;
5467: data <= 32'Hffffffeb;
5468: data <= 32'Hffffffed;
5469: data <= 32'Hffffffef;
5470: data <= 32'Hfffffff3;
5471: data <= 32'Hfffffff4;
5472: data <= 32'Hfffffff2;
5473: data <= 32'Hfffffff2;
5474: data <= 32'Hfffffff3;
5475: data <= 32'Hfffffff2;
5476: data <= 32'Hfffffff2;
5477: data <= 32'Hfffffff0;
5478: data <= 32'Hfffffff2;
5479: data <= 32'Hffffffef;
5480: data <= 32'Hffffffef;
5481: data <= 32'Hffffffee;
5482: data <= 32'Hffffffea;
5483: data <= 32'Hffffffe1;
5484: data <= 32'Hffffffdf;
5485: data <= 32'Hffffffde;
5486: data <= 32'Hffffffe3;
5487: data <= 32'Hffffffe6;
5488: data <= 32'Hffffffe2;
5489: data <= 32'Hffffffe2;
5490: data <= 32'Hffffffe7;
5491: data <= 32'Hffffffec;
5492: data <= 32'Hfffffff2;
5493: data <= 32'Hfffffff7;
5494: data <= 32'Hfffffff7;
5495: data <= 32'Hfffffff7;
5496: data <= 32'Hfffffff6;
5497: data <= 32'Hfffffffb;
5498: data <= 32'Hfffffff7;
5499: data <= 32'Hfffffff3;
5500: data <= 32'Hfffffff6;
5501: data <= 32'Hfffffff4;
5502: data <= 32'Hfffffffc;
5503: data <= 32'H00000000;
5504: data <= 32'H00000004;
5505: data <= 32'H00000006;
5506: data <= 32'H00000007;
5507: data <= 32'H00000004;
5508: data <= 32'H00000005;
5509: data <= 32'H00000009;
5510: data <= 32'H00000005;
5511: data <= 32'H00000004;
5512: data <= 32'H00000009;
5513: data <= 32'H00000005;
5514: data <= 32'H00000006;
5515: data <= 32'H00000005;
5516: data <= 32'H00000003;
5517: data <= 32'H00000007;
5518: data <= 32'H00000006;
5519: data <= 32'H00000004;
5520: data <= 32'H00000004;
5521: data <= 32'H00000005;
5522: data <= 32'H00000000;
5523: data <= 32'Hfffffff8;
5524: data <= 32'Hfffffff4;
5525: data <= 32'Hfffffff2;
5526: data <= 32'Hfffffff3;
5527: data <= 32'Hfffffffe;
5528: data <= 32'H00000005;
5529: data <= 32'H00000006;
5530: data <= 32'H00000004;
5531: data <= 32'H00000002;
5532: data <= 32'Hfffffffe;
5533: data <= 32'Hfffffff9;
5534: data <= 32'Hfffffff1;
5535: data <= 32'Hffffffef;
5536: data <= 32'Hfffffff2;
5537: data <= 32'Hfffffff5;
5538: data <= 32'Hfffffff7;
5539: data <= 32'Hfffffffc;
5540: data <= 32'Hfffffff9;
5541: data <= 32'H00000000;
5542: data <= 32'H00000006;
5543: data <= 32'H0000000a;
5544: data <= 32'H00000008;
5545: data <= 32'H00000004;
5546: data <= 32'Hfffffffd;
5547: data <= 32'Hfffffffa;
5548: data <= 32'Hfffffffb;
5549: data <= 32'Hfffffffb;
5550: data <= 32'Hfffffff8;
5551: data <= 32'Hfffffff8;
5552: data <= 32'Hfffffffe;
5553: data <= 32'H00000009;
5554: data <= 32'H0000000e;
5555: data <= 32'H00000007;
5556: data <= 32'Hfffffffa;
5557: data <= 32'Hfffffff8;
5558: data <= 32'Hfffffff6;
5559: data <= 32'Hfffffff6;
5560: data <= 32'Hffffffef;
5561: data <= 32'Hffffffea;
5562: data <= 32'Hffffffe2;
5563: data <= 32'Hffffffdc;
5564: data <= 32'Hffffffde;
5565: data <= 32'Hffffffe2;
5566: data <= 32'Hffffffeb;
5567: data <= 32'Hfffffff0;
5568: data <= 32'Hfffffff3;
5569: data <= 32'Hfffffff2;
5570: data <= 32'Hfffffff1;
5571: data <= 32'Hffffffed;
5572: data <= 32'Hffffffe8;
5573: data <= 32'Hffffffe6;
5574: data <= 32'Hffffffde;
5575: data <= 32'Hffffffd9;
5576: data <= 32'Hffffffd6;
5577: data <= 32'Hffffffcf;
5578: data <= 32'Hffffffd0;
5579: data <= 32'Hffffffd6;
5580: data <= 32'Hffffffd8;
5581: data <= 32'Hffffffd6;
5582: data <= 32'Hffffffd9;
5583: data <= 32'Hffffffda;
5584: data <= 32'Hffffffd7;
5585: data <= 32'Hffffffdb;
5586: data <= 32'Hffffffdc;
5587: data <= 32'Hffffffde;
5588: data <= 32'Hffffffe1;
5589: data <= 32'Hffffffde;
5590: data <= 32'Hffffffdd;
5591: data <= 32'Hffffffde;
5592: data <= 32'Hffffffe0;
5593: data <= 32'Hffffffe2;
5594: data <= 32'Hffffffe7;
5595: data <= 32'Hffffffeb;
5596: data <= 32'Hffffffea;
5597: data <= 32'Hffffffee;
5598: data <= 32'Hfffffff6;
5599: data <= 32'Hfffffff6;
5600: data <= 32'Hfffffff6;
5601: data <= 32'Hfffffff4;
5602: data <= 32'Hfffffff6;
5603: data <= 32'Hfffffff3;
5604: data <= 32'Hfffffff4;
5605: data <= 32'Hfffffff3;
5606: data <= 32'Hfffffff4;
5607: data <= 32'Hfffffff4;
5608: data <= 32'Hffffffee;
5609: data <= 32'Hffffffe8;
5610: data <= 32'Hffffffea;
5611: data <= 32'Hffffffe9;
5612: data <= 32'Hffffffeb;
5613: data <= 32'Hffffffe6;
5614: data <= 32'Hffffffe6;
5615: data <= 32'Hffffffe1;
5616: data <= 32'Hffffffdb;
5617: data <= 32'Hffffffdf;
5618: data <= 32'Hffffffe7;
5619: data <= 32'Hffffffea;
5620: data <= 32'Hfffffff1;
5621: data <= 32'Hfffffff9;
5622: data <= 32'Hfffffff7;
5623: data <= 32'Hfffffffb;
5624: data <= 32'Hfffffffb;
5625: data <= 32'Hfffffff6;
5626: data <= 32'Hfffffff6;
5627: data <= 32'Hfffffff4;
5628: data <= 32'Hfffffffa;
5629: data <= 32'Hffffffff;
5630: data <= 32'H00000001;
5631: data <= 32'H00000000;
5632: data <= 32'H00000007;
5633: data <= 32'H00000006;
5634: data <= 32'H00000005;
5635: data <= 32'H00000008;
5636: data <= 32'H00000006;
5637: data <= 32'H00000006;
5638: data <= 32'H00000007;
5639: data <= 32'H00000009;
5640: data <= 32'H00000005;
5641: data <= 32'H00000007;
5642: data <= 32'H00000005;
5643: data <= 32'H00000004;
5644: data <= 32'H00000005;
5645: data <= 32'H00000003;
5646: data <= 32'H00000004;
5647: data <= 32'H00000007;
5648: data <= 32'H00000002;
5649: data <= 32'H00000004;
5650: data <= 32'H00000003;
5651: data <= 32'Hfffffffd;
5652: data <= 32'Hfffffff7;
5653: data <= 32'Hfffffff0;
5654: data <= 32'Hffffffef;
5655: data <= 32'Hfffffff0;
5656: data <= 32'Hfffffffa;
5657: data <= 32'H00000003;
5658: data <= 32'H00000004;
5659: data <= 32'H00000001;
5660: data <= 32'H00000003;
5661: data <= 32'Hfffffffa;
5662: data <= 32'Hfffffff8;
5663: data <= 32'Hfffffff1;
5664: data <= 32'Hffffffed;
5665: data <= 32'Hfffffff1;
5666: data <= 32'Hffffffef;
5667: data <= 32'Hfffffff5;
5668: data <= 32'Hfffffffb;
5669: data <= 32'Hfffffffd;
5670: data <= 32'H00000001;
5671: data <= 32'H00000005;
5672: data <= 32'H0000000a;
5673: data <= 32'H0000000a;
5674: data <= 32'H00000003;
5675: data <= 32'Hfffffffc;
5676: data <= 32'Hfffffffd;
5677: data <= 32'Hfffffffd;
5678: data <= 32'Hfffffffd;
5679: data <= 32'Hfffffff9;
5680: data <= 32'Hfffffffa;
5681: data <= 32'H00000000;
5682: data <= 32'H00000007;
5683: data <= 32'H0000000e;
5684: data <= 32'H0000000a;
5685: data <= 32'H00000000;
5686: data <= 32'Hfffffff8;
5687: data <= 32'Hfffffff4;
5688: data <= 32'Hffffffee;
5689: data <= 32'Hffffffed;
5690: data <= 32'Hffffffe5;
5691: data <= 32'Hffffffe2;
5692: data <= 32'Hffffffe0;
5693: data <= 32'Hffffffe0;
5694: data <= 32'Hffffffe4;
5695: data <= 32'Hffffffea;
5696: data <= 32'Hfffffff1;
5697: data <= 32'Hfffffff3;
5698: data <= 32'Hfffffff2;
5699: data <= 32'Hfffffff0;
5700: data <= 32'Hffffffec;
5701: data <= 32'Hffffffe3;
5702: data <= 32'Hffffffe1;
5703: data <= 32'Hffffffdd;
5704: data <= 32'Hffffffd1;
5705: data <= 32'Hffffffd2;
5706: data <= 32'Hffffffd2;
5707: data <= 32'Hffffffd0;
5708: data <= 32'Hffffffd1;
5709: data <= 32'Hffffffd6;
5710: data <= 32'Hffffffd7;
5711: data <= 32'Hffffffd9;
5712: data <= 32'Hffffffda;
5713: data <= 32'Hffffffdd;
5714: data <= 32'Hffffffe1;
5715: data <= 32'Hffffffe2;
5716: data <= 32'Hffffffe1;
5717: data <= 32'Hffffffe1;
5718: data <= 32'Hffffffdf;
5719: data <= 32'Hffffffde;
5720: data <= 32'Hffffffde;
5721: data <= 32'Hffffffe3;
5722: data <= 32'Hffffffe7;
5723: data <= 32'Hffffffea;
5724: data <= 32'Hffffffef;
5725: data <= 32'Hfffffff2;
5726: data <= 32'Hfffffffa;
5727: data <= 32'Hfffffffe;
5728: data <= 32'Hfffffffe;
5729: data <= 32'Hfffffffc;
5730: data <= 32'Hffffffff;
5731: data <= 32'Hfffffffd;
5732: data <= 32'Hfffffffa;
5733: data <= 32'Hfffffff8;
5734: data <= 32'Hfffffff5;
5735: data <= 32'Hfffffff3;
5736: data <= 32'Hfffffff3;
5737: data <= 32'Hfffffff5;
5738: data <= 32'Hfffffff8;
5739: data <= 32'Hfffffff8;
5740: data <= 32'Hffffffed;
5741: data <= 32'Hffffffe3;
5742: data <= 32'Hffffffde;
5743: data <= 32'Hffffffdb;
5744: data <= 32'Hffffffdf;
5745: data <= 32'Hffffffe5;
5746: data <= 32'Hffffffea;
5747: data <= 32'Hffffffee;
5748: data <= 32'Hfffffff5;
5749: data <= 32'Hfffffff8;
5750: data <= 32'Hfffffffb;
5751: data <= 32'Hfffffff7;
5752: data <= 32'Hfffffff6;
5753: data <= 32'Hfffffff8;
5754: data <= 32'Hfffffffc;
5755: data <= 32'Hfffffffc;
5756: data <= 32'Hffffffff;
5757: data <= 32'Hfffffffb;
5758: data <= 32'H00000000;
5759: data <= 32'H00000001;
5760: data <= 32'Hffffffff;
5761: data <= 32'H00000005;
5762: data <= 32'H00000007;
5763: data <= 32'H00000008;
5764: data <= 32'H00000005;
5765: data <= 32'H00000008;
5766: data <= 32'H00000004;
5767: data <= 32'H00000007;
5768: data <= 32'H00000005;
5769: data <= 32'H00000006;
5770: data <= 32'H00000004;
5771: data <= 32'H00000004;
5772: data <= 32'H00000005;
5773: data <= 32'H00000002;
5774: data <= 32'H00000003;
5775: data <= 32'H00000005;
5776: data <= 32'H00000006;
5777: data <= 32'H00000003;
5778: data <= 32'H00000003;
5779: data <= 32'H00000001;
5780: data <= 32'Hfffffffe;
5781: data <= 32'Hfffffffb;
5782: data <= 32'Hfffffff3;
5783: data <= 32'Hfffffff0;
5784: data <= 32'Hfffffff2;
5785: data <= 32'Hfffffff7;
5786: data <= 32'H00000001;
5787: data <= 32'H00000004;
5788: data <= 32'H00000002;
5789: data <= 32'H00000004;
5790: data <= 32'Hfffffffe;
5791: data <= 32'Hfffffff7;
5792: data <= 32'Hfffffff6;
5793: data <= 32'Hfffffff1;
5794: data <= 32'Hffffffee;
5795: data <= 32'Hfffffff1;
5796: data <= 32'Hfffffff5;
5797: data <= 32'Hfffffffb;
5798: data <= 32'H00000000;
5799: data <= 32'Hffffffff;
5800: data <= 32'H00000006;
5801: data <= 32'H00000009;
5802: data <= 32'H00000007;
5803: data <= 32'H00000006;
5804: data <= 32'H00000002;
5805: data <= 32'Hfffffffc;
5806: data <= 32'Hffffffff;
5807: data <= 32'Hfffffffd;
5808: data <= 32'Hfffffff9;
5809: data <= 32'Hfffffffb;
5810: data <= 32'Hffffffff;
5811: data <= 32'H00000003;
5812: data <= 32'H0000000b;
5813: data <= 32'H0000000a;
5814: data <= 32'H00000005;
5815: data <= 32'Hfffffffe;
5816: data <= 32'Hfffffff1;
5817: data <= 32'Hfffffff1;
5818: data <= 32'Hffffffec;
5819: data <= 32'Hffffffee;
5820: data <= 32'Hffffffe8;
5821: data <= 32'Hffffffe7;
5822: data <= 32'Hffffffe6;
5823: data <= 32'Hffffffea;
5824: data <= 32'Hffffffed;
5825: data <= 32'Hfffffff1;
5826: data <= 32'Hfffffff4;
5827: data <= 32'Hfffffff4;
5828: data <= 32'Hfffffff1;
5829: data <= 32'Hffffffed;
5830: data <= 32'Hffffffe7;
5831: data <= 32'Hffffffe1;
5832: data <= 32'Hffffffdc;
5833: data <= 32'Hffffffd8;
5834: data <= 32'Hffffffd7;
5835: data <= 32'Hffffffd6;
5836: data <= 32'Hffffffd6;
5837: data <= 32'Hffffffdc;
5838: data <= 32'Hffffffdf;
5839: data <= 32'Hffffffe0;
5840: data <= 32'Hffffffe1;
5841: data <= 32'Hffffffe7;
5842: data <= 32'Hffffffe8;
5843: data <= 32'Hffffffe9;
5844: data <= 32'Hffffffe7;
5845: data <= 32'Hffffffe6;
5846: data <= 32'Hffffffe4;
5847: data <= 32'Hffffffe3;
5848: data <= 32'Hffffffe3;
5849: data <= 32'Hffffffe4;
5850: data <= 32'Hffffffea;
5851: data <= 32'Hffffffef;
5852: data <= 32'Hfffffff3;
5853: data <= 32'Hfffffff9;
5854: data <= 32'H00000000;
5855: data <= 32'H00000006;
5856: data <= 32'H00000007;
5857: data <= 32'H00000006;
5858: data <= 32'H00000007;
5859: data <= 32'H00000004;
5860: data <= 32'H00000002;
5861: data <= 32'Hfffffffe;
5862: data <= 32'Hfffffffe;
5863: data <= 32'H00000001;
5864: data <= 32'H00000002;
5865: data <= 32'Hffffffff;
5866: data <= 32'H00000001;
5867: data <= 32'Hfffffffb;
5868: data <= 32'Hffffffef;
5869: data <= 32'Hffffffe4;
5870: data <= 32'Hffffffe4;
5871: data <= 32'Hffffffe5;
5872: data <= 32'Hffffffea;
5873: data <= 32'Hffffffed;
5874: data <= 32'Hfffffff1;
5875: data <= 32'Hfffffff2;
5876: data <= 32'Hfffffff6;
5877: data <= 32'Hfffffff9;
5878: data <= 32'Hfffffff7;
5879: data <= 32'Hfffffff9;
5880: data <= 32'Hfffffffe;
5881: data <= 32'Hfffffffd;
5882: data <= 32'H00000002;
5883: data <= 32'Hffffffff;
5884: data <= 32'Hfffffffe;
5885: data <= 32'H00000000;
5886: data <= 32'H00000003;
5887: data <= 32'Hffffffff;
5888: data <= 32'H00000008;
5889: data <= 32'H00000007;
5890: data <= 32'H00000005;
5891: data <= 32'H00000006;
5892: data <= 32'H00000006;
5893: data <= 32'H00000007;
5894: data <= 32'H00000006;
5895: data <= 32'H00000006;
5896: data <= 32'H00000006;
5897: data <= 32'H00000004;
5898: data <= 32'H00000005;
5899: data <= 32'H00000005;
5900: data <= 32'H00000004;
5901: data <= 32'H00000005;
5902: data <= 32'H00000004;
5903: data <= 32'H00000001;
5904: data <= 32'H00000006;
5905: data <= 32'H00000005;
5906: data <= 32'H00000000;
5907: data <= 32'H00000003;
5908: data <= 32'H00000003;
5909: data <= 32'H00000000;
5910: data <= 32'Hfffffffe;
5911: data <= 32'Hfffffff9;
5912: data <= 32'Hfffffff2;
5913: data <= 32'Hfffffff4;
5914: data <= 32'Hfffffff3;
5915: data <= 32'Hfffffff9;
5916: data <= 32'H00000000;
5917: data <= 32'H00000002;
5918: data <= 32'H00000000;
5919: data <= 32'H00000000;
5920: data <= 32'Hfffffffb;
5921: data <= 32'Hfffffff6;
5922: data <= 32'Hfffffff1;
5923: data <= 32'Hffffffef;
5924: data <= 32'Hfffffff1;
5925: data <= 32'Hfffffff2;
5926: data <= 32'Hfffffff9;
5927: data <= 32'Hfffffffe;
5928: data <= 32'H00000002;
5929: data <= 32'H00000006;
5930: data <= 32'H00000008;
5931: data <= 32'H00000009;
5932: data <= 32'H0000000a;
5933: data <= 32'H00000004;
5934: data <= 32'H00000000;
5935: data <= 32'Hfffffffd;
5936: data <= 32'Hfffffffd;
5937: data <= 32'Hfffffffc;
5938: data <= 32'Hfffffff9;
5939: data <= 32'Hfffffffa;
5940: data <= 32'Hfffffffd;
5941: data <= 32'H00000007;
5942: data <= 32'H0000000d;
5943: data <= 32'H00000008;
5944: data <= 32'Hfffffffe;
5945: data <= 32'Hfffffff5;
5946: data <= 32'Hffffffef;
5947: data <= 32'Hffffffef;
5948: data <= 32'Hffffffee;
5949: data <= 32'Hffffffec;
5950: data <= 32'Hffffffec;
5951: data <= 32'Hffffffeb;
5952: data <= 32'Hffffffe8;
5953: data <= 32'Hffffffeb;
5954: data <= 32'Hffffffef;
5955: data <= 32'Hfffffff1;
5956: data <= 32'Hfffffff1;
5957: data <= 32'Hfffffff0;
5958: data <= 32'Hffffffee;
5959: data <= 32'Hffffffe7;
5960: data <= 32'Hffffffdf;
5961: data <= 32'Hffffffe0;
5962: data <= 32'Hffffffde;
5963: data <= 32'Hffffffdc;
5964: data <= 32'Hffffffde;
5965: data <= 32'Hffffffe4;
5966: data <= 32'Hffffffe6;
5967: data <= 32'Hffffffe6;
5968: data <= 32'Hffffffe9;
5969: data <= 32'Hffffffeb;
5970: data <= 32'Hffffffe9;
5971: data <= 32'Hffffffed;
5972: data <= 32'Hffffffee;
5973: data <= 32'Hffffffed;
5974: data <= 32'Hffffffe9;
5975: data <= 32'Hffffffe6;
5976: data <= 32'Hffffffe5;
5977: data <= 32'Hffffffe7;
5978: data <= 32'Hffffffe9;
5979: data <= 32'Hffffffef;
5980: data <= 32'Hfffffff5;
5981: data <= 32'Hfffffffd;
5982: data <= 32'H00000003;
5983: data <= 32'H00000006;
5984: data <= 32'H0000000b;
5985: data <= 32'H00000008;
5986: data <= 32'H00000007;
5987: data <= 32'H00000005;
5988: data <= 32'H00000006;
5989: data <= 32'H00000006;
5990: data <= 32'H00000009;
5991: data <= 32'H00000007;
5992: data <= 32'H00000007;
5993: data <= 32'H00000002;
5994: data <= 32'Hfffffffc;
5995: data <= 32'Hfffffff9;
5996: data <= 32'Hfffffff5;
5997: data <= 32'Hfffffff0;
5998: data <= 32'Hfffffff1;
5999: data <= 32'Hfffffff0;
6000: data <= 32'Hffffffed;
6001: data <= 32'Hfffffff2;
6002: data <= 32'Hfffffff7;
6003: data <= 32'Hfffffff2;
6004: data <= 32'Hfffffff6;
6005: data <= 32'Hfffffff6;
6006: data <= 32'Hfffffff7;
6007: data <= 32'Hfffffffc;
6008: data <= 32'Hfffffffe;
6009: data <= 32'Hfffffffb;
6010: data <= 32'Hffffffff;
6011: data <= 32'H00000000;
6012: data <= 32'H00000002;
6013: data <= 32'H00000005;
6014: data <= 32'H00000005;
6015: data <= 32'H00000007;
6016: data <= 32'H00000001;
6017: data <= 32'H00000007;
6018: data <= 32'H00000008;
6019: data <= 32'H00000008;
6020: data <= 32'H00000007;
6021: data <= 32'H00000007;
6022: data <= 32'H00000008;
6023: data <= 32'H00000007;
6024: data <= 32'H00000007;
6025: data <= 32'H00000009;
6026: data <= 32'H00000007;
6027: data <= 32'H00000006;
6028: data <= 32'H00000008;
6029: data <= 32'H00000006;
6030: data <= 32'H00000007;
6031: data <= 32'H00000006;
6032: data <= 32'H00000007;
6033: data <= 32'H00000006;
6034: data <= 32'H00000008;
6035: data <= 32'H00000007;
6036: data <= 32'H00000009;
6037: data <= 32'H00000008;
6038: data <= 32'H00000004;
6039: data <= 32'H00000006;
6040: data <= 32'H00000001;
6041: data <= 32'Hfffffffb;
6042: data <= 32'Hfffffff6;
6043: data <= 32'Hfffffff5;
6044: data <= 32'Hfffffff4;
6045: data <= 32'Hffffffff;
6046: data <= 32'H00000004;
6047: data <= 32'H00000007;
6048: data <= 32'H00000005;
6049: data <= 32'Hfffffffd;
6050: data <= 32'Hfffffff8;
6051: data <= 32'Hfffffff4;
6052: data <= 32'Hfffffff2;
6053: data <= 32'Hfffffff0;
6054: data <= 32'Hfffffff2;
6055: data <= 32'Hfffffff5;
6056: data <= 32'Hfffffffc;
6057: data <= 32'H00000006;
6058: data <= 32'H00000005;
6059: data <= 32'H00000009;
6060: data <= 32'H0000000b;
6061: data <= 32'H0000000b;
6062: data <= 32'H00000007;
6063: data <= 32'H00000005;
6064: data <= 32'Hffffffff;
6065: data <= 32'H00000002;
6066: data <= 32'H00000000;
6067: data <= 32'Hfffffffb;
6068: data <= 32'Hfffffffc;
6069: data <= 32'Hfffffffd;
6070: data <= 32'H00000006;
6071: data <= 32'H0000000d;
6072: data <= 32'H0000000c;
6073: data <= 32'H00000002;
6074: data <= 32'Hfffffff9;
6075: data <= 32'Hfffffff1;
6076: data <= 32'Hfffffff1;
6077: data <= 32'Hfffffff4;
6078: data <= 32'Hffffffee;
6079: data <= 32'Hffffffef;
6080: data <= 32'Hffffffed;
6081: data <= 32'Hffffffeb;
6082: data <= 32'Hffffffed;
6083: data <= 32'Hffffffec;
6084: data <= 32'Hfffffff0;
6085: data <= 32'Hfffffff1;
6086: data <= 32'Hfffffff1;
6087: data <= 32'Hffffffeb;
6088: data <= 32'Hffffffe9;
6089: data <= 32'Hffffffe8;
6090: data <= 32'Hffffffe6;
6091: data <= 32'Hffffffe3;
6092: data <= 32'Hffffffe8;
6093: data <= 32'Hffffffed;
6094: data <= 32'Hffffffec;
6095: data <= 32'Hffffffec;
6096: data <= 32'Hffffffee;
6097: data <= 32'Hfffffff0;
6098: data <= 32'Hfffffff0;
6099: data <= 32'Hfffffff1;
6100: data <= 32'Hfffffff0;
6101: data <= 32'Hfffffff5;
6102: data <= 32'Hfffffff0;
6103: data <= 32'Hffffffee;
6104: data <= 32'Hffffffee;
6105: data <= 32'Hffffffed;
6106: data <= 32'Hffffffef;
6107: data <= 32'Hfffffff3;
6108: data <= 32'Hfffffff9;
6109: data <= 32'Hfffffffd;
6110: data <= 32'H00000003;
6111: data <= 32'H00000008;
6112: data <= 32'H00000009;
6113: data <= 32'H0000000a;
6114: data <= 32'H0000000c;
6115: data <= 32'H0000000b;
6116: data <= 32'H0000000e;
6117: data <= 32'H0000000c;
6118: data <= 32'H0000000c;
6119: data <= 32'H00000008;
6120: data <= 32'H00000006;
6121: data <= 32'Hfffffffd;
6122: data <= 32'H00000002;
6123: data <= 32'Hfffffffe;
6124: data <= 32'H00000001;
6125: data <= 32'Hffffffff;
6126: data <= 32'Hfffffffe;
6127: data <= 32'Hfffffffd;
6128: data <= 32'Hfffffffd;
6129: data <= 32'Hfffffff8;
6130: data <= 32'Hfffffff3;
6131: data <= 32'Hfffffff1;
6132: data <= 32'Hfffffff4;
6133: data <= 32'Hfffffff5;
6134: data <= 32'Hfffffff5;
6135: data <= 32'Hfffffff3;
6136: data <= 32'Hfffffff4;
6137: data <= 32'Hfffffff8;
6138: data <= 32'H00000000;
6139: data <= 32'H00000004;
6140: data <= 32'H00000009;
6141: data <= 32'H00000009;
6142: data <= 32'H00000009;
6143: data <= 32'H00000004;
6144: data <= 32'H00000000;
6145: data <= 32'H00000009;
6146: data <= 32'H0000000a;
6147: data <= 32'H0000000a;
6148: data <= 32'H0000000a;
6149: data <= 32'H0000000a;
6150: data <= 32'H0000000a;
6151: data <= 32'H00000009;
6152: data <= 32'H0000000e;
6153: data <= 32'H00000009;
6154: data <= 32'H0000000a;
6155: data <= 32'H0000000b;
6156: data <= 32'H00000009;
6157: data <= 32'H0000000a;
6158: data <= 32'H0000000b;
6159: data <= 32'H00000008;
6160: data <= 32'H0000000b;
6161: data <= 32'H0000000c;
6162: data <= 32'H0000000d;
6163: data <= 32'H0000000c;
6164: data <= 32'H0000000b;
6165: data <= 32'H0000000b;
6166: data <= 32'H00000009;
6167: data <= 32'H0000000c;
6168: data <= 32'H0000000b;
6169: data <= 32'H00000007;
6170: data <= 32'H00000002;
6171: data <= 32'Hfffffffd;
6172: data <= 32'Hfffffff8;
6173: data <= 32'Hfffffff6;
6174: data <= 32'Hfffffffc;
6175: data <= 32'H00000004;
6176: data <= 32'H00000007;
6177: data <= 32'H00000008;
6178: data <= 32'H00000004;
6179: data <= 32'Hffffffff;
6180: data <= 32'Hfffffffb;
6181: data <= 32'Hfffffff5;
6182: data <= 32'Hfffffff2;
6183: data <= 32'Hfffffff4;
6184: data <= 32'Hfffffff3;
6185: data <= 32'Hfffffffa;
6186: data <= 32'Hffffffff;
6187: data <= 32'H00000001;
6188: data <= 32'H00000006;
6189: data <= 32'H00000008;
6190: data <= 32'H00000007;
6191: data <= 32'H00000007;
6192: data <= 32'H00000003;
6193: data <= 32'H00000000;
6194: data <= 32'H00000005;
6195: data <= 32'H00000001;
6196: data <= 32'Hffffffff;
6197: data <= 32'Hfffffffa;
6198: data <= 32'Hfffffffd;
6199: data <= 32'H00000001;
6200: data <= 32'H00000009;
6201: data <= 32'H0000000e;
6202: data <= 32'H00000009;
6203: data <= 32'H00000002;
6204: data <= 32'Hfffffffc;
6205: data <= 32'Hfffffffc;
6206: data <= 32'Hfffffff6;
6207: data <= 32'Hfffffff6;
6208: data <= 32'Hfffffff4;
6209: data <= 32'Hfffffff2;
6210: data <= 32'Hfffffff0;
6211: data <= 32'Hffffffef;
6212: data <= 32'Hfffffff1;
6213: data <= 32'Hfffffff2;
6214: data <= 32'Hfffffff4;
6215: data <= 32'Hfffffff0;
6216: data <= 32'Hfffffff4;
6217: data <= 32'Hfffffffa;
6218: data <= 32'Hfffffff1;
6219: data <= 32'Hfffffff0;
6220: data <= 32'Hfffffff2;
6221: data <= 32'Hfffffff4;
6222: data <= 32'Hfffffff6;
6223: data <= 32'Hfffffff4;
6224: data <= 32'Hfffffff7;
6225: data <= 32'Hfffffffb;
6226: data <= 32'Hfffffff8;
6227: data <= 32'Hfffffff9;
6228: data <= 32'Hfffffffa;
6229: data <= 32'Hfffffffb;
6230: data <= 32'Hfffffffa;
6231: data <= 32'Hfffffff8;
6232: data <= 32'Hfffffff8;
6233: data <= 32'Hfffffff9;
6234: data <= 32'Hfffffffa;
6235: data <= 32'H00000000;
6236: data <= 32'H00000003;
6237: data <= 32'H00000006;
6238: data <= 32'H0000000c;
6239: data <= 32'H00000012;
6240: data <= 32'H00000013;
6241: data <= 32'H00000017;
6242: data <= 32'H0000001a;
6243: data <= 32'H00000015;
6244: data <= 32'H00000014;
6245: data <= 32'H0000000e;
6246: data <= 32'H0000000c;
6247: data <= 32'H0000000b;
6248: data <= 32'H00000009;
6249: data <= 32'H00000008;
6250: data <= 32'H0000000b;
6251: data <= 32'H0000000b;
6252: data <= 32'H0000000e;
6253: data <= 32'H0000000d;
6254: data <= 32'H0000000c;
6255: data <= 32'H00000002;
6256: data <= 32'Hfffffff8;
6257: data <= 32'Hfffffff7;
6258: data <= 32'Hfffffff0;
6259: data <= 32'Hfffffff1;
6260: data <= 32'Hfffffff3;
6261: data <= 32'Hffffffed;
6262: data <= 32'Hffffffec;
6263: data <= 32'Hffffffee;
6264: data <= 32'Hfffffff1;
6265: data <= 32'Hfffffff6;
6266: data <= 32'H00000002;
6267: data <= 32'H00000007;
6268: data <= 32'H0000000a;
6269: data <= 32'H00000009;
6270: data <= 32'H00000005;
6271: data <= 32'H00000002;
6272: data <= 32'H00000000;
6273: data <= 32'H00000012;
6274: data <= 32'H00000011;
6275: data <= 32'H00000013;
6276: data <= 32'H00000015;
6277: data <= 32'H00000012;
6278: data <= 32'H00000012;
6279: data <= 32'H00000015;
6280: data <= 32'H00000012;
6281: data <= 32'H00000014;
6282: data <= 32'H00000014;
6283: data <= 32'H00000013;
6284: data <= 32'H00000014;
6285: data <= 32'H00000011;
6286: data <= 32'H00000010;
6287: data <= 32'H00000013;
6288: data <= 32'H00000015;
6289: data <= 32'H00000012;
6290: data <= 32'H00000013;
6291: data <= 32'H00000012;
6292: data <= 32'H00000013;
6293: data <= 32'H00000013;
6294: data <= 32'H00000017;
6295: data <= 32'H00000015;
6296: data <= 32'H00000015;
6297: data <= 32'H00000014;
6298: data <= 32'H00000011;
6299: data <= 32'H00000010;
6300: data <= 32'H0000000b;
6301: data <= 32'H00000006;
6302: data <= 32'Hfffffffe;
6303: data <= 32'Hfffffffd;
6304: data <= 32'Hffffffff;
6305: data <= 32'H00000006;
6306: data <= 32'H0000000b;
6307: data <= 32'H0000000c;
6308: data <= 32'H0000000f;
6309: data <= 32'H00000007;
6310: data <= 32'H00000000;
6311: data <= 32'Hfffffffe;
6312: data <= 32'Hfffffffa;
6313: data <= 32'Hfffffff9;
6314: data <= 32'Hfffffffb;
6315: data <= 32'Hfffffffd;
6316: data <= 32'H00000002;
6317: data <= 32'H0000000a;
6318: data <= 32'H0000000c;
6319: data <= 32'H00000011;
6320: data <= 32'H0000000e;
6321: data <= 32'H00000009;
6322: data <= 32'H0000000b;
6323: data <= 32'H00000004;
6324: data <= 32'H00000007;
6325: data <= 32'H00000008;
6326: data <= 32'H00000005;
6327: data <= 32'H00000006;
6328: data <= 32'H00000006;
6329: data <= 32'H0000000d;
6330: data <= 32'H00000010;
6331: data <= 32'H00000015;
6332: data <= 32'H0000000f;
6333: data <= 32'H0000000b;
6334: data <= 32'H00000007;
6335: data <= 32'H00000003;
6336: data <= 32'Hffffffff;
6337: data <= 32'H00000000;
6338: data <= 32'Hffffffff;
6339: data <= 32'Hfffffffc;
6340: data <= 32'Hfffffffe;
6341: data <= 32'H00000001;
6342: data <= 32'H00000001;
6343: data <= 32'H00000003;
6344: data <= 32'H00000002;
6345: data <= 32'H00000006;
6346: data <= 32'H00000003;
6347: data <= 32'Hfffffffd;
6348: data <= 32'Hfffffffb;
6349: data <= 32'H00000004;
6350: data <= 32'Hfffffffd;
6351: data <= 32'H00000004;
6352: data <= 32'H00000007;
6353: data <= 32'H00000006;
6354: data <= 32'H00000006;
6355: data <= 32'H00000008;
6356: data <= 32'H00000006;
6357: data <= 32'H0000000a;
6358: data <= 32'H0000000b;
6359: data <= 32'H0000000a;
6360: data <= 32'H00000009;
6361: data <= 32'H0000000b;
6362: data <= 32'H0000000c;
6363: data <= 32'H00000011;
6364: data <= 32'H00000017;
6365: data <= 32'H0000001b;
6366: data <= 32'H00000020;
6367: data <= 32'H00000026;
6368: data <= 32'H00000024;
6369: data <= 32'H00000025;
6370: data <= 32'H00000023;
6371: data <= 32'H0000001d;
6372: data <= 32'H00000018;
6373: data <= 32'H00000014;
6374: data <= 32'H00000013;
6375: data <= 32'H00000012;
6376: data <= 32'H00000011;
6377: data <= 32'H00000014;
6378: data <= 32'H00000018;
6379: data <= 32'H00000015;
6380: data <= 32'H00000012;
6381: data <= 32'H0000000c;
6382: data <= 32'H00000007;
6383: data <= 32'H00000003;
6384: data <= 32'Hfffffffe;
6385: data <= 32'Hfffffffb;
6386: data <= 32'Hfffffff1;
6387: data <= 32'Hfffffff8;
6388: data <= 32'Hfffffff3;
6389: data <= 32'Hfffffff4;
6390: data <= 32'Hfffffff6;
6391: data <= 32'Hfffffff8;
6392: data <= 32'Hfffffffd;
6393: data <= 32'H00000000;
6394: data <= 32'Hfffffffe;
6395: data <= 32'H00000000;
6396: data <= 32'Hfffffffe;
6397: data <= 32'Hfffffffe;
6398: data <= 32'H00000006;
6399: data <= 32'H00000006;
6400: data <= 32'H00000007;
6401: data <= 32'H0000000e;
6402: data <= 32'H0000000f;
6403: data <= 32'H00000010;
6404: data <= 32'H00000010;
6405: data <= 32'H00000012;
6406: data <= 32'H0000000e;
6407: data <= 32'H00000011;
6408: data <= 32'H0000000e;
6409: data <= 32'H0000000e;
6410: data <= 32'H00000012;
6411: data <= 32'H00000011;
6412: data <= 32'H0000000d;
6413: data <= 32'H00000010;
6414: data <= 32'H0000000e;
6415: data <= 32'H0000000f;
6416: data <= 32'H00000012;
6417: data <= 32'H00000011;
6418: data <= 32'H0000000e;
6419: data <= 32'H00000010;
6420: data <= 32'H00000010;
6421: data <= 32'H00000012;
6422: data <= 32'H00000011;
6423: data <= 32'H00000012;
6424: data <= 32'H00000012;
6425: data <= 32'H00000012;
6426: data <= 32'H00000011;
6427: data <= 32'H00000011;
6428: data <= 32'H00000012;
6429: data <= 32'H0000000e;
6430: data <= 32'H0000000b;
6431: data <= 32'H00000002;
6432: data <= 32'Hfffffffe;
6433: data <= 32'Hfffffffa;
6434: data <= 32'H00000000;
6435: data <= 32'H00000002;
6436: data <= 32'H0000000c;
6437: data <= 32'H00000010;
6438: data <= 32'H0000000e;
6439: data <= 32'H0000000c;
6440: data <= 32'H00000009;
6441: data <= 32'H00000001;
6442: data <= 32'H00000001;
6443: data <= 32'Hfffffffb;
6444: data <= 32'Hfffffffa;
6445: data <= 32'Hffffffff;
6446: data <= 32'H00000001;
6447: data <= 32'H00000008;
6448: data <= 32'H0000000e;
6449: data <= 32'H0000000f;
6450: data <= 32'H00000010;
6451: data <= 32'H0000000f;
6452: data <= 32'H00000008;
6453: data <= 32'H0000000a;
6454: data <= 32'H0000000a;
6455: data <= 32'H00000009;
6456: data <= 32'H00000006;
6457: data <= 32'H00000006;
6458: data <= 32'H00000007;
6459: data <= 32'H00000007;
6460: data <= 32'H0000000d;
6461: data <= 32'H00000010;
6462: data <= 32'H00000011;
6463: data <= 32'H00000010;
6464: data <= 32'H0000000a;
6465: data <= 32'H00000009;
6466: data <= 32'H00000008;
6467: data <= 32'H00000007;
6468: data <= 32'H00000003;
6469: data <= 32'H00000007;
6470: data <= 32'H00000006;
6471: data <= 32'H00000008;
6472: data <= 32'H00000004;
6473: data <= 32'H00000008;
6474: data <= 32'H00000004;
6475: data <= 32'H00000002;
6476: data <= 32'Hfffffff8;
6477: data <= 32'Hfffffff8;
6478: data <= 32'Hfffffffd;
6479: data <= 32'Hfffffffd;
6480: data <= 32'Hffffffff;
6481: data <= 32'H00000005;
6482: data <= 32'H00000006;
6483: data <= 32'H00000007;
6484: data <= 32'H0000000b;
6485: data <= 32'H0000000d;
6486: data <= 32'H0000000c;
6487: data <= 32'H00000010;
6488: data <= 32'H0000000f;
6489: data <= 32'H00000013;
6490: data <= 32'H00000016;
6491: data <= 32'H0000001a;
6492: data <= 32'H0000001f;
6493: data <= 32'H00000021;
6494: data <= 32'H00000025;
6495: data <= 32'H00000024;
6496: data <= 32'H00000023;
6497: data <= 32'H0000001e;
6498: data <= 32'H0000001a;
6499: data <= 32'H00000017;
6500: data <= 32'H00000017;
6501: data <= 32'H00000014;
6502: data <= 32'H0000001a;
6503: data <= 32'H00000017;
6504: data <= 32'H00000018;
6505: data <= 32'H00000015;
6506: data <= 32'H00000011;
6507: data <= 32'H00000010;
6508: data <= 32'H00000009;
6509: data <= 32'H00000006;
6510: data <= 32'Hffffffff;
6511: data <= 32'Hfffffffc;
6512: data <= 32'Hfffffff9;
6513: data <= 32'Hfffffffc;
6514: data <= 32'Hfffffff8;
6515: data <= 32'Hfffffffb;
6516: data <= 32'Hfffffff9;
6517: data <= 32'Hfffffff8;
6518: data <= 32'Hfffffff6;
6519: data <= 32'Hfffffff7;
6520: data <= 32'Hfffffff4;
6521: data <= 32'Hffffffec;
6522: data <= 32'Hffffffee;
6523: data <= 32'Hffffffed;
6524: data <= 32'Hffffffef;
6525: data <= 32'Hfffffffa;
6526: data <= 32'Hfffffffa;
6527: data <= 32'Hfffffffb;
6528: data <= 32'H00000000;
6529: data <= 32'H0000000a;
6530: data <= 32'H00000005;
6531: data <= 32'H00000005;
6532: data <= 32'H00000005;
6533: data <= 32'H00000007;
6534: data <= 32'H00000006;
6535: data <= 32'H00000008;
6536: data <= 32'H00000006;
6537: data <= 32'H00000005;
6538: data <= 32'H00000005;
6539: data <= 32'H00000005;
6540: data <= 32'H00000002;
6541: data <= 32'H00000003;
6542: data <= 32'H00000002;
6543: data <= 32'H00000003;
6544: data <= 32'H00000007;
6545: data <= 32'H00000005;
6546: data <= 32'H00000005;
6547: data <= 32'H0000000c;
6548: data <= 32'H0000000c;
6549: data <= 32'H0000000b;
6550: data <= 32'H0000000d;
6551: data <= 32'H0000000a;
6552: data <= 32'H0000000c;
6553: data <= 32'H00000010;
6554: data <= 32'H00000008;
6555: data <= 32'H00000008;
6556: data <= 32'H0000000c;
6557: data <= 32'H00000007;
6558: data <= 32'H00000007;
6559: data <= 32'H0000000a;
6560: data <= 32'H00000004;
6561: data <= 32'Hfffffffb;
6562: data <= 32'Hfffffffb;
6563: data <= 32'Hfffffff4;
6564: data <= 32'Hfffffff7;
6565: data <= 32'Hfffffffb;
6566: data <= 32'Hfffffffe;
6567: data <= 32'H00000005;
6568: data <= 32'H00000006;
6569: data <= 32'H00000000;
6570: data <= 32'H0000000a;
6571: data <= 32'H00000001;
6572: data <= 32'Hfffffffa;
6573: data <= 32'Hfffffffd;
6574: data <= 32'Hffffffef;
6575: data <= 32'Hfffffff5;
6576: data <= 32'Hfffffffe;
6577: data <= 32'H00000003;
6578: data <= 32'H00000008;
6579: data <= 32'H0000000e;
6580: data <= 32'H0000000d;
6581: data <= 32'H00000007;
6582: data <= 32'H00000006;
6583: data <= 32'H00000004;
6584: data <= 32'H00000004;
6585: data <= 32'H00000001;
6586: data <= 32'Hffffffff;
6587: data <= 32'Hfffffffb;
6588: data <= 32'Hfffffffe;
6589: data <= 32'Hfffffffd;
6590: data <= 32'H00000000;
6591: data <= 32'H00000007;
6592: data <= 32'H00000007;
6593: data <= 32'H00000008;
6594: data <= 32'H0000000c;
6595: data <= 32'H0000000b;
6596: data <= 32'H0000000c;
6597: data <= 32'H0000000d;
6598: data <= 32'H0000000b;
6599: data <= 32'H0000000b;
6600: data <= 32'H00000007;
6601: data <= 32'H0000000a;
6602: data <= 32'H00000006;
6603: data <= 32'H00000003;
6604: data <= 32'Hfffffffc;
6605: data <= 32'Hfffffffa;
6606: data <= 32'Hfffffff9;
6607: data <= 32'Hfffffffc;
6608: data <= 32'Hffffffff;
6609: data <= 32'H00000002;
6610: data <= 32'H00000004;
6611: data <= 32'H00000009;
6612: data <= 32'H0000000a;
6613: data <= 32'H0000000d;
6614: data <= 32'H0000000d;
6615: data <= 32'H00000012;
6616: data <= 32'H00000012;
6617: data <= 32'H00000013;
6618: data <= 32'H00000016;
6619: data <= 32'H00000019;
6620: data <= 32'H00000017;
6621: data <= 32'H0000001b;
6622: data <= 32'H00000018;
6623: data <= 32'H00000014;
6624: data <= 32'H00000016;
6625: data <= 32'H00000013;
6626: data <= 32'H00000011;
6627: data <= 32'H00000018;
6628: data <= 32'H00000018;
6629: data <= 32'H00000015;
6630: data <= 32'H00000017;
6631: data <= 32'H0000000f;
6632: data <= 32'H0000000b;
6633: data <= 32'H00000006;
6634: data <= 32'H00000000;
6635: data <= 32'Hffffffff;
6636: data <= 32'Hfffffffb;
6637: data <= 32'Hfffffffb;
6638: data <= 32'Hfffffff9;
6639: data <= 32'Hfffffffd;
6640: data <= 32'Hffffffff;
6641: data <= 32'Hfffffffe;
6642: data <= 32'Hfffffffb;
6643: data <= 32'Hffffffff;
6644: data <= 32'Hfffffffa;
6645: data <= 32'Hfffffff3;
6646: data <= 32'Hfffffff2;
6647: data <= 32'Hffffffec;
6648: data <= 32'Hffffffe3;
6649: data <= 32'Hffffffe4;
6650: data <= 32'Hffffffe5;
6651: data <= 32'Hffffffe4;
6652: data <= 32'Hffffffec;
6653: data <= 32'Hfffffff0;
6654: data <= 32'Hfffffff2;
6655: data <= 32'Hfffffff0;
6656: data <= 32'Hfffffff0;
6657: data <= 32'H0000000b;
6658: data <= 32'H0000000d;
6659: data <= 32'H0000000e;
6660: data <= 32'H0000000d;
6661: data <= 32'H0000000e;
6662: data <= 32'H00000011;
6663: data <= 32'H0000000a;
6664: data <= 32'H0000000b;
6665: data <= 32'H0000000e;
6666: data <= 32'H00000009;
6667: data <= 32'H0000000b;
6668: data <= 32'H0000000c;
6669: data <= 32'H0000000c;
6670: data <= 32'H0000000b;
6671: data <= 32'H0000000a;
6672: data <= 32'H0000000b;
6673: data <= 32'H0000000d;
6674: data <= 32'H00000010;
6675: data <= 32'H0000000e;
6676: data <= 32'H00000012;
6677: data <= 32'H00000013;
6678: data <= 32'H0000000c;
6679: data <= 32'H00000011;
6680: data <= 32'H00000014;
6681: data <= 32'H0000000c;
6682: data <= 32'H00000010;
6683: data <= 32'H00000011;
6684: data <= 32'H0000000a;
6685: data <= 32'H0000000f;
6686: data <= 32'H00000010;
6687: data <= 32'H00000007;
6688: data <= 32'H0000000c;
6689: data <= 32'H0000000c;
6690: data <= 32'H00000008;
6691: data <= 32'H00000005;
6692: data <= 32'H00000000;
6693: data <= 32'Hfffffffb;
6694: data <= 32'Hfffffffb;
6695: data <= 32'Hfffffffc;
6696: data <= 32'Hfffffffc;
6697: data <= 32'Hfffffffd;
6698: data <= 32'H00000006;
6699: data <= 32'H00000007;
6700: data <= 32'Hfffffff8;
6701: data <= 32'H00000002;
6702: data <= 32'Hfffffff0;
6703: data <= 32'Hffffffe5;
6704: data <= 32'Hffffffee;
6705: data <= 32'Hffffffea;
6706: data <= 32'Hffffffef;
6707: data <= 32'Hfffffffe;
6708: data <= 32'H00000004;
6709: data <= 32'H00000006;
6710: data <= 32'H00000008;
6711: data <= 32'H00000007;
6712: data <= 32'H00000007;
6713: data <= 32'H00000000;
6714: data <= 32'H00000008;
6715: data <= 32'H0000000a;
6716: data <= 32'H00000006;
6717: data <= 32'H00000008;
6718: data <= 32'H00000004;
6719: data <= 32'H00000003;
6720: data <= 32'H00000004;
6721: data <= 32'H00000006;
6722: data <= 32'H00000011;
6723: data <= 32'H00000016;
6724: data <= 32'H00000018;
6725: data <= 32'H00000019;
6726: data <= 32'H00000021;
6727: data <= 32'H0000001a;
6728: data <= 32'H00000017;
6729: data <= 32'H00000015;
6730: data <= 32'H0000000b;
6731: data <= 32'H0000000c;
6732: data <= 32'H00000003;
6733: data <= 32'Hffffffff;
6734: data <= 32'Hfffffffa;
6735: data <= 32'Hfffffff9;
6736: data <= 32'Hffffffff;
6737: data <= 32'Hffffffff;
6738: data <= 32'Hffffffff;
6739: data <= 32'H00000009;
6740: data <= 32'H00000007;
6741: data <= 32'H0000000f;
6742: data <= 32'H0000000d;
6743: data <= 32'H00000010;
6744: data <= 32'H00000010;
6745: data <= 32'H0000000e;
6746: data <= 32'H0000000d;
6747: data <= 32'H00000011;
6748: data <= 32'H0000000e;
6749: data <= 32'H0000000f;
6750: data <= 32'H00000010;
6751: data <= 32'H00000012;
6752: data <= 32'H00000015;
6753: data <= 32'H00000018;
6754: data <= 32'H0000001a;
6755: data <= 32'H0000001d;
6756: data <= 32'H0000001c;
6757: data <= 32'H00000011;
6758: data <= 32'H0000000f;
6759: data <= 32'H0000000d;
6760: data <= 32'H00000003;
6761: data <= 32'H00000002;
6762: data <= 32'H00000000;
6763: data <= 32'H00000001;
6764: data <= 32'H00000004;
6765: data <= 32'H0000000e;
6766: data <= 32'H0000000d;
6767: data <= 32'H0000000e;
6768: data <= 32'H0000000e;
6769: data <= 32'H0000000e;
6770: data <= 32'H0000000c;
6771: data <= 32'H00000012;
6772: data <= 32'H0000000c;
6773: data <= 32'H00000002;
6774: data <= 32'Hfffffffc;
6775: data <= 32'Hfffffffb;
6776: data <= 32'Hfffffff4;
6777: data <= 32'Hfffffff4;
6778: data <= 32'Hfffffff9;
6779: data <= 32'Hfffffff3;
6780: data <= 32'Hfffffff6;
6781: data <= 32'H00000000;
6782: data <= 32'Hfffffffd;
6783: data <= 32'Hffffffff;
6784: data <= 32'H00000004;
6785: data <= 32'H00000009;
6786: data <= 32'H0000000b;
6787: data <= 32'H0000000c;
6788: data <= 32'H0000000e;
6789: data <= 32'H0000000b;
6790: data <= 32'H0000000e;
6791: data <= 32'H0000000d;
6792: data <= 32'H0000000a;
6793: data <= 32'H0000000e;
6794: data <= 32'H0000000e;
6795: data <= 32'H0000000e;
6796: data <= 32'H0000000b;
6797: data <= 32'H0000000f;
6798: data <= 32'H0000000e;
6799: data <= 32'H0000000b;
6800: data <= 32'H0000000e;
6801: data <= 32'H0000000e;
6802: data <= 32'H0000000d;
6803: data <= 32'H00000011;
6804: data <= 32'H00000012;
6805: data <= 32'H0000000d;
6806: data <= 32'H00000010;
6807: data <= 32'H00000010;
6808: data <= 32'H0000000c;
6809: data <= 32'H0000000e;
6810: data <= 32'H0000000f;
6811: data <= 32'H0000000d;
6812: data <= 32'H0000000d;
6813: data <= 32'H00000011;
6814: data <= 32'H0000000e;
6815: data <= 32'H0000000d;
6816: data <= 32'H0000000d;
6817: data <= 32'H0000000d;
6818: data <= 32'H0000000d;
6819: data <= 32'H0000000c;
6820: data <= 32'H00000010;
6821: data <= 32'H0000000e;
6822: data <= 32'H00000007;
6823: data <= 32'H00000003;
6824: data <= 32'Hfffffffc;
6825: data <= 32'Hfffffffa;
6826: data <= 32'Hfffffffe;
6827: data <= 32'H00000000;
6828: data <= 32'Hfffffffe;
6829: data <= 32'H00000005;
6830: data <= 32'H00000007;
6831: data <= 32'Hfffffffe;
6832: data <= 32'H00000003;
6833: data <= 32'Hfffffffa;
6834: data <= 32'Hffffffef;
6835: data <= 32'Hfffffff2;
6836: data <= 32'Hffffffec;
6837: data <= 32'Hffffffec;
6838: data <= 32'Hfffffff7;
6839: data <= 32'Hfffffffc;
6840: data <= 32'Hfffffffb;
6841: data <= 32'Hffffffff;
6842: data <= 32'H00000003;
6843: data <= 32'H00000003;
6844: data <= 32'H00000004;
6845: data <= 32'H00000008;
6846: data <= 32'H0000000c;
6847: data <= 32'H00000009;
6848: data <= 32'H0000000a;
6849: data <= 32'H0000000b;
6850: data <= 32'H0000000c;
6851: data <= 32'H0000000f;
6852: data <= 32'H00000010;
6853: data <= 32'H00000014;
6854: data <= 32'H0000001c;
6855: data <= 32'H0000001a;
6856: data <= 32'H0000001d;
6857: data <= 32'H00000019;
6858: data <= 32'H00000017;
6859: data <= 32'H00000013;
6860: data <= 32'H0000000b;
6861: data <= 32'H00000006;
6862: data <= 32'H00000002;
6863: data <= 32'Hfffffff8;
6864: data <= 32'Hfffffff8;
6865: data <= 32'Hfffffff8;
6866: data <= 32'Hfffffff3;
6867: data <= 32'Hfffffff7;
6868: data <= 32'Hfffffff9;
6869: data <= 32'Hfffffffe;
6870: data <= 32'Hfffffffd;
6871: data <= 32'H00000002;
6872: data <= 32'H00000004;
6873: data <= 32'H00000003;
6874: data <= 32'H0000000d;
6875: data <= 32'H00000010;
6876: data <= 32'H00000012;
6877: data <= 32'H00000019;
6878: data <= 32'H0000001b;
6879: data <= 32'H0000001d;
6880: data <= 32'H00000021;
6881: data <= 32'H0000001b;
6882: data <= 32'H00000016;
6883: data <= 32'H00000014;
6884: data <= 32'H0000000d;
6885: data <= 32'H00000007;
6886: data <= 32'H0000000c;
6887: data <= 32'H0000000d;
6888: data <= 32'H00000008;
6889: data <= 32'H0000000e;
6890: data <= 32'H0000000b;
6891: data <= 32'H0000000f;
6892: data <= 32'H00000014;
6893: data <= 32'H00000019;
6894: data <= 32'H0000001b;
6895: data <= 32'H00000017;
6896: data <= 32'H00000016;
6897: data <= 32'H00000016;
6898: data <= 32'H0000001a;
6899: data <= 32'H0000001e;
6900: data <= 32'H00000019;
6901: data <= 32'H00000010;
6902: data <= 32'H00000003;
6903: data <= 32'Hfffffffb;
6904: data <= 32'Hfffffff5;
6905: data <= 32'Hfffffff6;
6906: data <= 32'Hfffffff9;
6907: data <= 32'Hfffffff8;
6908: data <= 32'Hfffffff9;
6909: data <= 32'Hfffffffe;
6910: data <= 32'Hfffffffe;
6911: data <= 32'H00000003;
6912: data <= 32'H00000008;
6913: data <= 32'H00000004;
6914: data <= 32'H00000005;
6915: data <= 32'H00000007;
6916: data <= 32'H00000006;
6917: data <= 32'H00000008;
6918: data <= 32'H00000008;
6919: data <= 32'H00000006;
6920: data <= 32'H00000006;
6921: data <= 32'H00000007;
6922: data <= 32'H00000008;
6923: data <= 32'H00000007;
6924: data <= 32'H00000008;
6925: data <= 32'H00000008;
6926: data <= 32'H00000006;
6927: data <= 32'H0000000d;
6928: data <= 32'H00000009;
6929: data <= 32'H00000005;
6930: data <= 32'H0000000c;
6931: data <= 32'H0000000b;
6932: data <= 32'H00000009;
6933: data <= 32'H0000000a;
6934: data <= 32'H0000000a;
6935: data <= 32'H00000009;
6936: data <= 32'H0000000c;
6937: data <= 32'H0000000a;
6938: data <= 32'H0000000a;
6939: data <= 32'H0000000a;
6940: data <= 32'H00000009;
6941: data <= 32'H00000009;
6942: data <= 32'H0000000a;
6943: data <= 32'H0000000c;
6944: data <= 32'H0000000a;
6945: data <= 32'H0000000a;
6946: data <= 32'H0000000b;
6947: data <= 32'H00000009;
6948: data <= 32'H00000006;
6949: data <= 32'H00000009;
6950: data <= 32'H0000000a;
6951: data <= 32'H0000000a;
6952: data <= 32'H0000000e;
6953: data <= 32'H00000008;
6954: data <= 32'H00000004;
6955: data <= 32'H00000001;
6956: data <= 32'Hfffffffa;
6957: data <= 32'Hfffffff7;
6958: data <= 32'Hfffffffd;
6959: data <= 32'Hfffffff9;
6960: data <= 32'Hfffffff9;
6961: data <= 32'H00000000;
6962: data <= 32'Hfffffff9;
6963: data <= 32'Hfffffffb;
6964: data <= 32'Hfffffffb;
6965: data <= 32'Hfffffff2;
6966: data <= 32'Hfffffff5;
6967: data <= 32'Hfffffff7;
6968: data <= 32'Hffffffef;
6969: data <= 32'Hfffffff3;
6970: data <= 32'Hfffffff7;
6971: data <= 32'Hfffffff4;
6972: data <= 32'Hffffffef;
6973: data <= 32'Hfffffff2;
6974: data <= 32'Hfffffff8;
6975: data <= 32'Hfffffff4;
6976: data <= 32'Hfffffffa;
6977: data <= 32'Hfffffffb;
6978: data <= 32'Hfffffff8;
6979: data <= 32'Hfffffffa;
6980: data <= 32'Hfffffffb;
6981: data <= 32'Hfffffffa;
6982: data <= 32'Hffffffff;
6983: data <= 32'H00000000;
6984: data <= 32'H00000006;
6985: data <= 32'H00000007;
6986: data <= 32'H0000000d;
6987: data <= 32'H0000000d;
6988: data <= 32'H0000000a;
6989: data <= 32'H00000006;
6990: data <= 32'H00000006;
6991: data <= 32'Hfffffff7;
6992: data <= 32'Hfffffff2;
6993: data <= 32'Hffffffed;
6994: data <= 32'Hffffffea;
6995: data <= 32'Hffffffe5;
6996: data <= 32'Hffffffea;
6997: data <= 32'Hffffffe8;
6998: data <= 32'Hfffffff1;
6999: data <= 32'Hfffffff2;
7000: data <= 32'Hfffffff6;
7001: data <= 32'Hfffffff9;
7002: data <= 32'H00000003;
7003: data <= 32'Hfffffffe;
7004: data <= 32'H00000003;
7005: data <= 32'H0000000a;
7006: data <= 32'H00000005;
7007: data <= 32'H00000002;
7008: data <= 32'H00000002;
7009: data <= 32'Hfffffff8;
7010: data <= 32'Hfffffff8;
7011: data <= 32'H00000000;
7012: data <= 32'Hfffffffc;
7013: data <= 32'H00000008;
7014: data <= 32'H0000000f;
7015: data <= 32'H00000010;
7016: data <= 32'H00000013;
7017: data <= 32'H00000015;
7018: data <= 32'H00000010;
7019: data <= 32'H00000013;
7020: data <= 32'H00000015;
7021: data <= 32'H00000014;
7022: data <= 32'H00000011;
7023: data <= 32'H00000014;
7024: data <= 32'H00000010;
7025: data <= 32'H00000011;
7026: data <= 32'H0000001c;
7027: data <= 32'H0000001c;
7028: data <= 32'H00000019;
7029: data <= 32'H00000018;
7030: data <= 32'H00000009;
7031: data <= 32'Hfffffff6;
7032: data <= 32'Hfffffff0;
7033: data <= 32'Hffffffee;
7034: data <= 32'Hffffffed;
7035: data <= 32'Hfffffff2;
7036: data <= 32'Hfffffff2;
7037: data <= 32'Hfffffff5;
7038: data <= 32'Hfffffff8;
7039: data <= 32'Hfffffffc;
7040: data <= 32'Hffffffff;
7041: data <= 32'H00000001;
7042: data <= 32'H00000001;
7043: data <= 32'H00000000;
7044: data <= 32'Hffffffff;
7045: data <= 32'H00000002;
7046: data <= 32'H00000003;
7047: data <= 32'H00000001;
7048: data <= 32'H00000004;
7049: data <= 32'H00000003;
7050: data <= 32'H00000001;
7051: data <= 32'H00000003;
7052: data <= 32'H00000002;
7053: data <= 32'H00000002;
7054: data <= 32'H00000004;
7055: data <= 32'H00000005;
7056: data <= 32'H00000003;
7057: data <= 32'H00000006;
7058: data <= 32'H00000003;
7059: data <= 32'H00000003;
7060: data <= 32'H00000005;
7061: data <= 32'H00000007;
7062: data <= 32'H00000003;
7063: data <= 32'H00000003;
7064: data <= 32'H00000006;
7065: data <= 32'H00000003;
7066: data <= 32'H00000004;
7067: data <= 32'H00000005;
7068: data <= 32'H00000004;
7069: data <= 32'Hffffffff;
7070: data <= 32'H00000003;
7071: data <= 32'H00000003;
7072: data <= 32'H00000002;
7073: data <= 32'H00000002;
7074: data <= 32'H00000006;
7075: data <= 32'H00000004;
7076: data <= 32'H00000001;
7077: data <= 32'H00000000;
7078: data <= 32'H00000002;
7079: data <= 32'H00000002;
7080: data <= 32'H00000004;
7081: data <= 32'H00000005;
7082: data <= 32'H00000005;
7083: data <= 32'H00000006;
7084: data <= 32'H00000005;
7085: data <= 32'H00000001;
7086: data <= 32'Hfffffffe;
7087: data <= 32'Hfffffff9;
7088: data <= 32'Hfffffff9;
7089: data <= 32'Hfffffff8;
7090: data <= 32'Hffffffee;
7091: data <= 32'Hffffffed;
7092: data <= 32'Hffffffee;
7093: data <= 32'Hffffffea;
7094: data <= 32'Hffffffeb;
7095: data <= 32'Hffffffef;
7096: data <= 32'Hffffffea;
7097: data <= 32'Hffffffef;
7098: data <= 32'Hfffffff4;
7099: data <= 32'Hfffffff5;
7100: data <= 32'Hfffffff5;
7101: data <= 32'Hfffffff8;
7102: data <= 32'Hfffffff7;
7103: data <= 32'Hfffffff6;
7104: data <= 32'Hfffffff9;
7105: data <= 32'Hfffffff6;
7106: data <= 32'Hfffffff6;
7107: data <= 32'Hfffffff5;
7108: data <= 32'Hffffffee;
7109: data <= 32'Hffffffea;
7110: data <= 32'Hffffffec;
7111: data <= 32'Hffffffea;
7112: data <= 32'Hffffffe9;
7113: data <= 32'Hffffffeb;
7114: data <= 32'Hfffffff0;
7115: data <= 32'Hfffffff1;
7116: data <= 32'Hfffffffc;
7117: data <= 32'Hfffffff2;
7118: data <= 32'H00000001;
7119: data <= 32'Hfffffffc;
7120: data <= 32'Hfffffff8;
7121: data <= 32'Hfffffff9;
7122: data <= 32'Hfffffffa;
7123: data <= 32'Hffffffed;
7124: data <= 32'Hfffffff9;
7125: data <= 32'Hffffffea;
7126: data <= 32'Hfffffff0;
7127: data <= 32'Hffffffef;
7128: data <= 32'Hfffffff0;
7129: data <= 32'Hffffffec;
7130: data <= 32'Hfffffff2;
7131: data <= 32'Hffffffe9;
7132: data <= 32'Hffffffeb;
7133: data <= 32'Hffffffee;
7134: data <= 32'Hffffffee;
7135: data <= 32'Hffffffec;
7136: data <= 32'Hfffffff5;
7137: data <= 32'Hfffffff8;
7138: data <= 32'Hfffffffb;
7139: data <= 32'H00000006;
7140: data <= 32'H00000006;
7141: data <= 32'H0000000f;
7142: data <= 32'H00000007;
7143: data <= 32'H00000005;
7144: data <= 32'H00000008;
7145: data <= 32'H00000001;
7146: data <= 32'Hfffffffa;
7147: data <= 32'H00000002;
7148: data <= 32'Hffffffff;
7149: data <= 32'H00000003;
7150: data <= 32'H00000006;
7151: data <= 32'H0000000c;
7152: data <= 32'H00000004;
7153: data <= 32'H00000009;
7154: data <= 32'H0000000a;
7155: data <= 32'H0000000b;
7156: data <= 32'H0000000e;
7157: data <= 32'H0000000c;
7158: data <= 32'H00000002;
7159: data <= 32'Hfffffff6;
7160: data <= 32'Hffffffeb;
7161: data <= 32'Hffffffea;
7162: data <= 32'Hfffffff0;
7163: data <= 32'Hfffffff3;
7164: data <= 32'Hfffffff4;
7165: data <= 32'Hfffffff7;
7166: data <= 32'Hfffffff7;
7167: data <= 32'Hfffffff7;
7168: data <= 32'Hfffffffd;
7169: data <= 32'Hffffffff;
7170: data <= 32'Hfffffffb;
7171: data <= 32'Hfffffffc;
7172: data <= 32'Hfffffffb;
7173: data <= 32'Hffffffff;
7174: data <= 32'Hfffffffd;
7175: data <= 32'H00000003;
7176: data <= 32'Hfffffffc;
7177: data <= 32'H00000000;
7178: data <= 32'Hfffffffe;
7179: data <= 32'Hfffffffe;
7180: data <= 32'Hfffffffc;
7181: data <= 32'H00000003;
7182: data <= 32'Hffffffff;
7183: data <= 32'H00000003;
7184: data <= 32'H00000000;
7185: data <= 32'H00000002;
7186: data <= 32'H00000001;
7187: data <= 32'H00000001;
7188: data <= 32'H00000004;
7189: data <= 32'H00000001;
7190: data <= 32'H00000002;
7191: data <= 32'H00000002;
7192: data <= 32'H00000002;
7193: data <= 32'H00000002;
7194: data <= 32'H00000004;
7195: data <= 32'H00000002;
7196: data <= 32'H00000002;
7197: data <= 32'Hffffffff;
7198: data <= 32'H00000003;
7199: data <= 32'Hffffffff;
7200: data <= 32'H00000003;
7201: data <= 32'Hfffffffd;
7202: data <= 32'H00000006;
7203: data <= 32'Hfffffffe;
7204: data <= 32'H00000003;
7205: data <= 32'H00000001;
7206: data <= 32'H00000004;
7207: data <= 32'H00000003;
7208: data <= 32'H00000003;
7209: data <= 32'H00000002;
7210: data <= 32'H00000005;
7211: data <= 32'H00000003;
7212: data <= 32'H00000003;
7213: data <= 32'H00000005;
7214: data <= 32'H00000003;
7215: data <= 32'H00000004;
7216: data <= 32'H00000002;
7217: data <= 32'H00000002;
7218: data <= 32'Hfffffffd;
7219: data <= 32'Hfffffffb;
7220: data <= 32'Hfffffff8;
7221: data <= 32'Hfffffffb;
7222: data <= 32'Hfffffff5;
7223: data <= 32'Hfffffff9;
7224: data <= 32'Hffffffee;
7225: data <= 32'Hfffffff0;
7226: data <= 32'Hffffffed;
7227: data <= 32'Hffffffed;
7228: data <= 32'Hffffffe5;
7229: data <= 32'Hffffffed;
7230: data <= 32'Hffffffe4;
7231: data <= 32'Hffffffe5;
7232: data <= 32'Hffffffeb;
7233: data <= 32'Hffffffe5;
7234: data <= 32'Hffffffe8;
7235: data <= 32'Hffffffea;
7236: data <= 32'Hffffffe8;
7237: data <= 32'Hffffffe7;
7238: data <= 32'Hffffffe9;
7239: data <= 32'Hffffffe6;
7240: data <= 32'Hffffffeb;
7241: data <= 32'Hffffffe1;
7242: data <= 32'Hffffffe5;
7243: data <= 32'Hffffffe3;
7244: data <= 32'Hffffffeb;
7245: data <= 32'Hffffffe2;
7246: data <= 32'Hffffffeb;
7247: data <= 32'Hffffffee;
7248: data <= 32'Hfffffff5;
7249: data <= 32'Hfffffff6;
7250: data <= 32'Hffffffff;
7251: data <= 32'Hfffffff6;
7252: data <= 32'H00000003;
7253: data <= 32'Hfffffffc;
7254: data <= 32'Hfffffffc;
7255: data <= 32'Hfffffff9;
7256: data <= 32'Hfffffffe;
7257: data <= 32'Hfffffff5;
7258: data <= 32'Hffffffff;
7259: data <= 32'H00000002;
7260: data <= 32'Hfffffffe;
7261: data <= 32'H00000004;
7262: data <= 32'H00000008;
7263: data <= 32'H00000005;
7264: data <= 32'H00000006;
7265: data <= 32'H00000009;
7266: data <= 32'H00000003;
7267: data <= 32'H00000001;
7268: data <= 32'Hfffffffc;
7269: data <= 32'Hffffffff;
7270: data <= 32'Hfffffff4;
7271: data <= 32'Hfffffffa;
7272: data <= 32'Hfffffffa;
7273: data <= 32'Hfffffff5;
7274: data <= 32'Hfffffff1;
7275: data <= 32'Hfffffff5;
7276: data <= 32'Hffffffef;
7277: data <= 32'Hfffffff6;
7278: data <= 32'Hfffffff0;
7279: data <= 32'Hfffffff6;
7280: data <= 32'Hfffffff2;
7281: data <= 32'Hfffffff6;
7282: data <= 32'Hfffffffc;
7283: data <= 32'H00000002;
7284: data <= 32'H00000005;
7285: data <= 32'H0000000b;
7286: data <= 32'H00000000;
7287: data <= 32'Hfffffff6;
7288: data <= 32'Hfffffff2;
7289: data <= 32'Hfffffff0;
7290: data <= 32'Hfffffff5;
7291: data <= 32'Hfffffff6;
7292: data <= 32'Hfffffffb;
7293: data <= 32'Hfffffffc;
7294: data <= 32'H00000003;
7295: data <= 32'H00000004;
7296: data <= 32'H0000000a;
7297: data <= 32'Hffffffec;
7298: data <= 32'Hffffffef;
7299: data <= 32'Hfffffff6;
7300: data <= 32'Hffffffed;
7301: data <= 32'Hfffffff4;
7302: data <= 32'Hfffffff4;
7303: data <= 32'Hfffffff3;
7304: data <= 32'Hfffffff4;
7305: data <= 32'Hfffffff7;
7306: data <= 32'Hfffffff0;
7307: data <= 32'Hfffffff7;
7308: data <= 32'Hfffffff3;
7309: data <= 32'Hfffffff6;
7310: data <= 32'Hfffffff5;
7311: data <= 32'Hfffffff8;
7312: data <= 32'Hfffffff6;
7313: data <= 32'Hfffffff8;
7314: data <= 32'Hfffffff9;
7315: data <= 32'Hfffffff8;
7316: data <= 32'Hfffffffb;
7317: data <= 32'Hfffffffa;
7318: data <= 32'Hfffffff9;
7319: data <= 32'Hfffffffb;
7320: data <= 32'Hfffffffc;
7321: data <= 32'Hfffffff7;
7322: data <= 32'Hfffffffb;
7323: data <= 32'Hfffffff8;
7324: data <= 32'Hfffffff8;
7325: data <= 32'Hfffffff8;
7326: data <= 32'Hfffffffa;
7327: data <= 32'Hfffffff5;
7328: data <= 32'Hfffffffe;
7329: data <= 32'Hfffffff7;
7330: data <= 32'Hfffffffc;
7331: data <= 32'Hfffffffa;
7332: data <= 32'Hfffffffc;
7333: data <= 32'Hfffffffa;
7334: data <= 32'Hfffffffd;
7335: data <= 32'Hfffffffc;
7336: data <= 32'Hfffffffb;
7337: data <= 32'Hfffffffd;
7338: data <= 32'Hfffffffc;
7339: data <= 32'Hfffffffd;
7340: data <= 32'Hfffffffe;
7341: data <= 32'Hfffffffc;
7342: data <= 32'H00000001;
7343: data <= 32'Hffffffff;
7344: data <= 32'H00000000;
7345: data <= 32'H00000001;
7346: data <= 32'Hfffffffe;
7347: data <= 32'Hffffffff;
7348: data <= 32'Hfffffffa;
7349: data <= 32'Hfffffffc;
7350: data <= 32'Hfffffff6;
7351: data <= 32'Hfffffff9;
7352: data <= 32'Hfffffff2;
7353: data <= 32'Hfffffff4;
7354: data <= 32'Hfffffff2;
7355: data <= 32'Hfffffff5;
7356: data <= 32'Hfffffff1;
7357: data <= 32'Hfffffff6;
7358: data <= 32'Hfffffff3;
7359: data <= 32'Hfffffff2;
7360: data <= 32'Hfffffff3;
7361: data <= 32'Hfffffff3;
7362: data <= 32'Hffffffeb;
7363: data <= 32'Hfffffff0;
7364: data <= 32'Hfffffff0;
7365: data <= 32'Hffffffec;
7366: data <= 32'Hfffffff5;
7367: data <= 32'Hfffffff1;
7368: data <= 32'Hfffffff5;
7369: data <= 32'Hfffffff4;
7370: data <= 32'Hfffffff5;
7371: data <= 32'Hfffffff6;
7372: data <= 32'H00000000;
7373: data <= 32'Hfffffff8;
7374: data <= 32'Hfffffffc;
7375: data <= 32'Hfffffffd;
7376: data <= 32'H00000002;
7377: data <= 32'Hffffffff;
7378: data <= 32'H00000004;
7379: data <= 32'H00000000;
7380: data <= 32'H00000001;
7381: data <= 32'Hfffffffb;
7382: data <= 32'H00000003;
7383: data <= 32'Hfffffffa;
7384: data <= 32'H00000001;
7385: data <= 32'H00000001;
7386: data <= 32'H00000005;
7387: data <= 32'H00000007;
7388: data <= 32'H00000003;
7389: data <= 32'Hfffffffe;
7390: data <= 32'Hfffffffc;
7391: data <= 32'Hfffffff9;
7392: data <= 32'Hfffffff3;
7393: data <= 32'Hfffffff7;
7394: data <= 32'Hfffffff1;
7395: data <= 32'Hffffffec;
7396: data <= 32'Hffffffea;
7397: data <= 32'Hffffffea;
7398: data <= 32'Hffffffe4;
7399: data <= 32'Hffffffe7;
7400: data <= 32'Hffffffe3;
7401: data <= 32'Hffffffe5;
7402: data <= 32'Hffffffdd;
7403: data <= 32'Hffffffde;
7404: data <= 32'Hffffffda;
7405: data <= 32'Hffffffe1;
7406: data <= 32'Hffffffd8;
7407: data <= 32'Hffffffe2;
7408: data <= 32'Hffffffe3;
7409: data <= 32'Hffffffe8;
7410: data <= 32'Hffffffed;
7411: data <= 32'Hfffffff1;
7412: data <= 32'Hfffffff3;
7413: data <= 32'Hfffffff5;
7414: data <= 32'Hfffffff1;
7415: data <= 32'Hffffffeb;
7416: data <= 32'Hffffffe9;
7417: data <= 32'Hffffffed;
7418: data <= 32'Hfffffff3;
7419: data <= 32'Hfffffff2;
7420: data <= 32'Hfffffffc;
7421: data <= 32'Hfffffffe;
7422: data <= 32'H00000001;
7423: data <= 32'H00000006;
7424: data <= 32'H00000010;
7425: data <= 32'Hfffffff3;
7426: data <= 32'Hfffffff6;
7427: data <= 32'Hfffffff3;
7428: data <= 32'Hfffffff6;
7429: data <= 32'Hfffffff5;
7430: data <= 32'Hfffffff7;
7431: data <= 32'Hfffffff9;
7432: data <= 32'Hfffffffb;
7433: data <= 32'Hfffffffa;
7434: data <= 32'Hfffffffc;
7435: data <= 32'Hfffffffb;
7436: data <= 32'Hfffffffb;
7437: data <= 32'Hfffffffe;
7438: data <= 32'Hfffffffc;
7439: data <= 32'Hfffffffe;
7440: data <= 32'Hffffffff;
7441: data <= 32'Hffffffff;
7442: data <= 32'Hfffffffd;
7443: data <= 32'H00000000;
7444: data <= 32'Hffffffff;
7445: data <= 32'Hfffffffc;
7446: data <= 32'Hfffffffd;
7447: data <= 32'Hfffffffe;
7448: data <= 32'Hfffffffd;
7449: data <= 32'Hfffffffe;
7450: data <= 32'Hfffffffd;
7451: data <= 32'Hffffffff;
7452: data <= 32'Hffffffff;
7453: data <= 32'Hfffffffe;
7454: data <= 32'Hfffffffc;
7455: data <= 32'Hfffffffe;
7456: data <= 32'H00000000;
7457: data <= 32'Hfffffffd;
7458: data <= 32'Hffffffff;
7459: data <= 32'H00000001;
7460: data <= 32'H00000002;
7461: data <= 32'H00000000;
7462: data <= 32'Hffffffff;
7463: data <= 32'H00000002;
7464: data <= 32'H00000001;
7465: data <= 32'Hfffffffe;
7466: data <= 32'H00000000;
7467: data <= 32'H00000002;
7468: data <= 32'H00000002;
7469: data <= 32'H00000003;
7470: data <= 32'H00000003;
7471: data <= 32'H00000006;
7472: data <= 32'H00000005;
7473: data <= 32'H00000005;
7474: data <= 32'H00000003;
7475: data <= 32'H00000001;
7476: data <= 32'H00000002;
7477: data <= 32'H00000004;
7478: data <= 32'Hfffffffe;
7479: data <= 32'H00000000;
7480: data <= 32'Hfffffffe;
7481: data <= 32'Hfffffffd;
7482: data <= 32'Hfffffffb;
7483: data <= 32'Hfffffff8;
7484: data <= 32'Hfffffff8;
7485: data <= 32'Hfffffff8;
7486: data <= 32'Hfffffff6;
7487: data <= 32'Hfffffff8;
7488: data <= 32'Hfffffffa;
7489: data <= 32'Hfffffff9;
7490: data <= 32'Hfffffff7;
7491: data <= 32'Hfffffff9;
7492: data <= 32'Hfffffff4;
7493: data <= 32'Hfffffffb;
7494: data <= 32'Hfffffffc;
7495: data <= 32'Hfffffffa;
7496: data <= 32'Hfffffffb;
7497: data <= 32'Hfffffffa;
7498: data <= 32'Hfffffff8;
7499: data <= 32'Hfffffff6;
7500: data <= 32'Hfffffff8;
7501: data <= 32'Hfffffff6;
7502: data <= 32'Hfffffff3;
7503: data <= 32'Hfffffff4;
7504: data <= 32'Hfffffff5;
7505: data <= 32'Hfffffff3;
7506: data <= 32'Hfffffff3;
7507: data <= 32'Hfffffff4;
7508: data <= 32'Hffffffed;
7509: data <= 32'Hffffffef;
7510: data <= 32'Hfffffff2;
7511: data <= 32'Hffffffee;
7512: data <= 32'Hfffffff6;
7513: data <= 32'Hfffffffb;
7514: data <= 32'Hfffffffb;
7515: data <= 32'Hfffffffd;
7516: data <= 32'Hfffffffc;
7517: data <= 32'Hfffffff4;
7518: data <= 32'Hfffffff2;
7519: data <= 32'Hffffffed;
7520: data <= 32'Hffffffed;
7521: data <= 32'Hffffffea;
7522: data <= 32'Hffffffe6;
7523: data <= 32'Hffffffe7;
7524: data <= 32'Hffffffe5;
7525: data <= 32'Hffffffe4;
7526: data <= 32'Hffffffe1;
7527: data <= 32'Hffffffe9;
7528: data <= 32'Hffffffe7;
7529: data <= 32'Hffffffe8;
7530: data <= 32'Hffffffea;
7531: data <= 32'Hffffffe3;
7532: data <= 32'Hffffffe7;
7533: data <= 32'Hffffffe7;
7534: data <= 32'Hffffffe6;
7535: data <= 32'Hffffffe7;
7536: data <= 32'Hffffffeb;
7537: data <= 32'Hfffffff0;
7538: data <= 32'Hffffffee;
7539: data <= 32'Hfffffff0;
7540: data <= 32'Hfffffff0;
7541: data <= 32'Hfffffff2;
7542: data <= 32'Hfffffff1;
7543: data <= 32'Hfffffff1;
7544: data <= 32'Hfffffff4;
7545: data <= 32'Hfffffffa;
7546: data <= 32'Hfffffffd;
7547: data <= 32'H00000004;
7548: data <= 32'H00000004;
7549: data <= 32'H00000009;
7550: data <= 32'H0000000c;
7551: data <= 32'H0000000f;
7552: data <= 32'H00000013;
7553: data <= 32'Hffffffec;
7554: data <= 32'Hffffffef;
7555: data <= 32'Hfffffff0;
7556: data <= 32'Hffffffef;
7557: data <= 32'Hffffffee;
7558: data <= 32'Hfffffff4;
7559: data <= 32'Hfffffff0;
7560: data <= 32'Hfffffff4;
7561: data <= 32'Hfffffff6;
7562: data <= 32'Hfffffff5;
7563: data <= 32'Hfffffff5;
7564: data <= 32'Hfffffff9;
7565: data <= 32'Hfffffff7;
7566: data <= 32'Hfffffffa;
7567: data <= 32'Hfffffffb;
7568: data <= 32'Hfffffff8;
7569: data <= 32'Hfffffffa;
7570: data <= 32'Hfffffffb;
7571: data <= 32'Hfffffff7;
7572: data <= 32'Hfffffff6;
7573: data <= 32'Hfffffffc;
7574: data <= 32'Hfffffff9;
7575: data <= 32'Hfffffff8;
7576: data <= 32'Hfffffffc;
7577: data <= 32'Hfffffff6;
7578: data <= 32'Hfffffffc;
7579: data <= 32'Hfffffffb;
7580: data <= 32'Hfffffff9;
7581: data <= 32'Hfffffff8;
7582: data <= 32'Hfffffff9;
7583: data <= 32'Hfffffffb;
7584: data <= 32'Hfffffff8;
7585: data <= 32'Hfffffffd;
7586: data <= 32'Hfffffffa;
7587: data <= 32'Hfffffffd;
7588: data <= 32'Hfffffffa;
7589: data <= 32'Hfffffffd;
7590: data <= 32'Hfffffffd;
7591: data <= 32'Hfffffffc;
7592: data <= 32'Hfffffffe;
7593: data <= 32'Hffffffff;
7594: data <= 32'Hfffffffd;
7595: data <= 32'H00000000;
7596: data <= 32'Hfffffffe;
7597: data <= 32'Hfffffffd;
7598: data <= 32'Hffffffff;
7599: data <= 32'Hffffffff;
7600: data <= 32'Hffffffff;
7601: data <= 32'H00000002;
7602: data <= 32'H00000001;
7603: data <= 32'Hfffffffa;
7604: data <= 32'Hfffffffd;
7605: data <= 32'H00000001;
7606: data <= 32'Hfffffffb;
7607: data <= 32'Hfffffffb;
7608: data <= 32'Hfffffffe;
7609: data <= 32'Hfffffffc;
7610: data <= 32'Hfffffff9;
7611: data <= 32'Hfffffffc;
7612: data <= 32'Hfffffffc;
7613: data <= 32'Hfffffff9;
7614: data <= 32'Hfffffffa;
7615: data <= 32'Hfffffff9;
7616: data <= 32'Hfffffff9;
7617: data <= 32'Hfffffff8;
7618: data <= 32'Hfffffff3;
7619: data <= 32'Hfffffff5;
7620: data <= 32'Hfffffff5;
7621: data <= 32'Hfffffff5;
7622: data <= 32'Hfffffff6;
7623: data <= 32'Hfffffff6;
7624: data <= 32'Hfffffff3;
7625: data <= 32'Hfffffff5;
7626: data <= 32'Hfffffff3;
7627: data <= 32'Hfffffff4;
7628: data <= 32'Hfffffff1;
7629: data <= 32'Hfffffff7;
7630: data <= 32'Hfffffff3;
7631: data <= 32'Hfffffff2;
7632: data <= 32'Hfffffff3;
7633: data <= 32'Hfffffff2;
7634: data <= 32'Hfffffff0;
7635: data <= 32'Hfffffff1;
7636: data <= 32'Hffffffee;
7637: data <= 32'Hfffffff1;
7638: data <= 32'Hfffffff3;
7639: data <= 32'Hfffffff7;
7640: data <= 32'Hfffffff9;
7641: data <= 32'H00000000;
7642: data <= 32'Hfffffffb;
7643: data <= 32'Hfffffffb;
7644: data <= 32'Hfffffffd;
7645: data <= 32'Hfffffff0;
7646: data <= 32'Hfffffff4;
7647: data <= 32'Hfffffff2;
7648: data <= 32'Hffffffec;
7649: data <= 32'Hffffffed;
7650: data <= 32'Hffffffee;
7651: data <= 32'Hffffffeb;
7652: data <= 32'Hffffffec;
7653: data <= 32'Hffffffec;
7654: data <= 32'Hffffffe5;
7655: data <= 32'Hffffffe8;
7656: data <= 32'Hffffffea;
7657: data <= 32'Hffffffeb;
7658: data <= 32'Hffffffeb;
7659: data <= 32'Hffffffec;
7660: data <= 32'Hffffffef;
7661: data <= 32'Hffffffec;
7662: data <= 32'Hffffffed;
7663: data <= 32'Hffffffe9;
7664: data <= 32'Hfffffff0;
7665: data <= 32'Hffffffeb;
7666: data <= 32'Hffffffee;
7667: data <= 32'Hffffffed;
7668: data <= 32'Hffffffec;
7669: data <= 32'Hffffffef;
7670: data <= 32'Hfffffff1;
7671: data <= 32'Hfffffff2;
7672: data <= 32'Hfffffff9;
7673: data <= 32'Hfffffffd;
7674: data <= 32'Hfffffffe;
7675: data <= 32'H00000007;
7676: data <= 32'H00000006;
7677: data <= 32'H00000009;
7678: data <= 32'H0000000b;
7679: data <= 32'H00000011;
7680: data <= 32'H0000000d;
7681: data <= 32'Hffffffe8;
7682: data <= 32'Hffffffe8;
7683: data <= 32'Hffffffe9;
7684: data <= 32'Hffffffed;
7685: data <= 32'Hffffffea;
7686: data <= 32'Hffffffea;
7687: data <= 32'Hfffffff0;
7688: data <= 32'Hffffffee;
7689: data <= 32'Hffffffed;
7690: data <= 32'Hfffffff1;
7691: data <= 32'Hffffffef;
7692: data <= 32'Hfffffff3;
7693: data <= 32'Hfffffff1;
7694: data <= 32'Hfffffff5;
7695: data <= 32'Hfffffff5;
7696: data <= 32'Hfffffff4;
7697: data <= 32'Hfffffff3;
7698: data <= 32'Hfffffff4;
7699: data <= 32'Hfffffff3;
7700: data <= 32'Hfffffff5;
7701: data <= 32'Hfffffff3;
7702: data <= 32'Hfffffff9;
7703: data <= 32'Hfffffff6;
7704: data <= 32'Hfffffff6;
7705: data <= 32'Hfffffff8;
7706: data <= 32'Hfffffff8;
7707: data <= 32'Hfffffff6;
7708: data <= 32'Hfffffff7;
7709: data <= 32'Hfffffff6;
7710: data <= 32'Hfffffff5;
7711: data <= 32'Hfffffff9;
7712: data <= 32'Hfffffff8;
7713: data <= 32'Hfffffffb;
7714: data <= 32'Hfffffff7;
7715: data <= 32'Hfffffffa;
7716: data <= 32'Hfffffff7;
7717: data <= 32'Hfffffffb;
7718: data <= 32'Hfffffffb;
7719: data <= 32'Hfffffffc;
7720: data <= 32'Hfffffffb;
7721: data <= 32'Hfffffffd;
7722: data <= 32'Hfffffffe;
7723: data <= 32'Hfffffffb;
7724: data <= 32'Hfffffffd;
7725: data <= 32'Hfffffffd;
7726: data <= 32'Hfffffffd;
7727: data <= 32'Hfffffffd;
7728: data <= 32'Hfffffffd;
7729: data <= 32'Hffffffff;
7730: data <= 32'Hffffffff;
7731: data <= 32'Hfffffffb;
7732: data <= 32'Hfffffffc;
7733: data <= 32'Hfffffffb;
7734: data <= 32'Hfffffffb;
7735: data <= 32'Hfffffffb;
7736: data <= 32'Hfffffffa;
7737: data <= 32'Hfffffffb;
7738: data <= 32'Hfffffff9;
7739: data <= 32'Hfffffffe;
7740: data <= 32'Hfffffffb;
7741: data <= 32'Hfffffffb;
7742: data <= 32'Hfffffffa;
7743: data <= 32'Hfffffff9;
7744: data <= 32'Hfffffff6;
7745: data <= 32'Hfffffff6;
7746: data <= 32'Hfffffff9;
7747: data <= 32'Hfffffff2;
7748: data <= 32'Hfffffff6;
7749: data <= 32'Hfffffff5;
7750: data <= 32'Hfffffff3;
7751: data <= 32'Hfffffff4;
7752: data <= 32'Hfffffff3;
7753: data <= 32'Hffffffef;
7754: data <= 32'Hfffffff2;
7755: data <= 32'Hfffffff2;
7756: data <= 32'Hffffffef;
7757: data <= 32'Hfffffff2;
7758: data <= 32'Hffffffed;
7759: data <= 32'Hffffffed;
7760: data <= 32'Hffffffec;
7761: data <= 32'Hffffffed;
7762: data <= 32'Hffffffea;
7763: data <= 32'Hffffffe8;
7764: data <= 32'Hffffffe9;
7765: data <= 32'Hffffffea;
7766: data <= 32'Hffffffee;
7767: data <= 32'Hfffffff5;
7768: data <= 32'Hfffffff5;
7769: data <= 32'Hfffffffa;
7770: data <= 32'Hfffffffb;
7771: data <= 32'Hfffffffa;
7772: data <= 32'Hfffffff4;
7773: data <= 32'Hfffffff2;
7774: data <= 32'Hfffffff1;
7775: data <= 32'Hfffffff3;
7776: data <= 32'Hfffffff2;
7777: data <= 32'Hfffffff3;
7778: data <= 32'Hfffffff1;
7779: data <= 32'Hfffffff3;
7780: data <= 32'Hffffffef;
7781: data <= 32'Hfffffff2;
7782: data <= 32'Hffffffed;
7783: data <= 32'Hffffffed;
7784: data <= 32'Hffffffed;
7785: data <= 32'Hfffffff0;
7786: data <= 32'Hffffffee;
7787: data <= 32'Hffffffef;
7788: data <= 32'Hfffffff6;
7789: data <= 32'Hffffffed;
7790: data <= 32'Hfffffff2;
7791: data <= 32'Hfffffff0;
7792: data <= 32'Hfffffff4;
7793: data <= 32'Hffffffef;
7794: data <= 32'Hffffffee;
7795: data <= 32'Hffffffef;
7796: data <= 32'Hfffffff0;
7797: data <= 32'Hfffffff0;
7798: data <= 32'Hfffffff6;
7799: data <= 32'Hfffffffa;
7800: data <= 32'Hfffffffc;
7801: data <= 32'H00000000;
7802: data <= 32'H00000000;
7803: data <= 32'H00000009;
7804: data <= 32'H00000006;
7805: data <= 32'H00000009;
7806: data <= 32'H00000009;
7807: data <= 32'H0000000b;
7808: data <= 32'H0000000b;
7809: data <= 32'Hffffffe9;
7810: data <= 32'Hffffffe4;
7811: data <= 32'Hffffffe6;
7812: data <= 32'Hffffffe7;
7813: data <= 32'Hffffffea;
7814: data <= 32'Hffffffe7;
7815: data <= 32'Hffffffed;
7816: data <= 32'Hffffffeb;
7817: data <= 32'Hffffffec;
7818: data <= 32'Hffffffee;
7819: data <= 32'Hffffffee;
7820: data <= 32'Hffffffef;
7821: data <= 32'Hfffffff0;
7822: data <= 32'Hfffffff0;
7823: data <= 32'Hfffffff2;
7824: data <= 32'Hfffffff3;
7825: data <= 32'Hfffffff1;
7826: data <= 32'Hfffffff1;
7827: data <= 32'Hfffffff4;
7828: data <= 32'Hfffffff4;
7829: data <= 32'Hfffffff4;
7830: data <= 32'Hfffffff4;
7831: data <= 32'Hfffffff6;
7832: data <= 32'Hfffffff7;
7833: data <= 32'Hfffffff7;
7834: data <= 32'Hfffffff7;
7835: data <= 32'Hfffffff3;
7836: data <= 32'Hfffffff7;
7837: data <= 32'Hfffffff5;
7838: data <= 32'Hfffffff5;
7839: data <= 32'Hfffffff7;
7840: data <= 32'Hfffffffa;
7841: data <= 32'Hfffffff8;
7842: data <= 32'Hfffffff7;
7843: data <= 32'Hfffffff8;
7844: data <= 32'Hfffffff9;
7845: data <= 32'Hfffffffa;
7846: data <= 32'Hfffffffd;
7847: data <= 32'Hfffffffc;
7848: data <= 32'Hfffffffc;
7849: data <= 32'Hfffffffd;
7850: data <= 32'Hfffffffd;
7851: data <= 32'Hfffffffc;
7852: data <= 32'Hfffffffe;
7853: data <= 32'Hfffffffe;
7854: data <= 32'Hffffffff;
7855: data <= 32'H00000000;
7856: data <= 32'Hffffffff;
7857: data <= 32'Hffffffff;
7858: data <= 32'H00000001;
7859: data <= 32'Hffffffff;
7860: data <= 32'Hfffffffc;
7861: data <= 32'Hffffffff;
7862: data <= 32'Hfffffffd;
7863: data <= 32'Hfffffffb;
7864: data <= 32'Hfffffffa;
7865: data <= 32'Hfffffff9;
7866: data <= 32'Hfffffffb;
7867: data <= 32'Hfffffffe;
7868: data <= 32'Hfffffffc;
7869: data <= 32'Hfffffffc;
7870: data <= 32'Hfffffffd;
7871: data <= 32'Hfffffffa;
7872: data <= 32'Hfffffff7;
7873: data <= 32'Hfffffffa;
7874: data <= 32'Hfffffffa;
7875: data <= 32'Hfffffff8;
7876: data <= 32'Hfffffff8;
7877: data <= 32'Hfffffff7;
7878: data <= 32'Hfffffff6;
7879: data <= 32'Hfffffff3;
7880: data <= 32'Hfffffff6;
7881: data <= 32'Hffffffef;
7882: data <= 32'Hfffffff3;
7883: data <= 32'Hfffffff3;
7884: data <= 32'Hfffffff1;
7885: data <= 32'Hfffffff2;
7886: data <= 32'Hfffffff0;
7887: data <= 32'Hffffffee;
7888: data <= 32'Hfffffff0;
7889: data <= 32'Hffffffec;
7890: data <= 32'Hffffffee;
7891: data <= 32'Hffffffea;
7892: data <= 32'Hffffffec;
7893: data <= 32'Hffffffeb;
7894: data <= 32'Hffffffee;
7895: data <= 32'Hfffffff3;
7896: data <= 32'Hfffffff4;
7897: data <= 32'Hfffffffa;
7898: data <= 32'H00000003;
7899: data <= 32'H00000004;
7900: data <= 32'H00000000;
7901: data <= 32'Hfffffffe;
7902: data <= 32'Hfffffffd;
7903: data <= 32'H00000000;
7904: data <= 32'Hffffffff;
7905: data <= 32'Hfffffffe;
7906: data <= 32'Hfffffffb;
7907: data <= 32'H00000000;
7908: data <= 32'Hfffffff8;
7909: data <= 32'Hfffffffa;
7910: data <= 32'Hfffffffc;
7911: data <= 32'Hfffffffa;
7912: data <= 32'Hfffffff7;
7913: data <= 32'Hfffffffa;
7914: data <= 32'Hfffffff7;
7915: data <= 32'Hfffffff6;
7916: data <= 32'Hfffffff7;
7917: data <= 32'Hfffffff6;
7918: data <= 32'Hfffffff2;
7919: data <= 32'Hfffffff3;
7920: data <= 32'Hfffffff3;
7921: data <= 32'Hfffffff2;
7922: data <= 32'Hfffffff1;
7923: data <= 32'Hfffffff3;
7924: data <= 32'Hfffffff3;
7925: data <= 32'Hfffffff6;
7926: data <= 32'Hfffffffb;
7927: data <= 32'Hfffffffb;
7928: data <= 32'H00000001;
7929: data <= 32'H00000001;
7930: data <= 32'H00000002;
7931: data <= 32'H00000006;
7932: data <= 32'H00000004;
7933: data <= 32'H00000006;
7934: data <= 32'H00000005;
7935: data <= 32'H00000009;
7936: data <= 32'H00000008;
7937: data <= 32'Hffffffed;
7938: data <= 32'Hffffffed;
7939: data <= 32'Hffffffee;
7940: data <= 32'Hffffffe8;
7941: data <= 32'Hffffffec;
7942: data <= 32'Hffffffeb;
7943: data <= 32'Hffffffec;
7944: data <= 32'Hffffffed;
7945: data <= 32'Hfffffff1;
7946: data <= 32'Hfffffff1;
7947: data <= 32'Hfffffff1;
7948: data <= 32'Hfffffff4;
7949: data <= 32'Hfffffff3;
7950: data <= 32'Hfffffff7;
7951: data <= 32'Hfffffff8;
7952: data <= 32'Hfffffff6;
7953: data <= 32'Hfffffffa;
7954: data <= 32'Hfffffff8;
7955: data <= 32'Hfffffff8;
7956: data <= 32'Hfffffff9;
7957: data <= 32'Hfffffff7;
7958: data <= 32'Hfffffff8;
7959: data <= 32'Hfffffff9;
7960: data <= 32'Hfffffffa;
7961: data <= 32'Hfffffff9;
7962: data <= 32'Hfffffff7;
7963: data <= 32'Hfffffff8;
7964: data <= 32'Hfffffffa;
7965: data <= 32'Hfffffffb;
7966: data <= 32'Hfffffffa;
7967: data <= 32'Hfffffffa;
7968: data <= 32'Hfffffffd;
7969: data <= 32'Hfffffff8;
7970: data <= 32'Hfffffff9;
7971: data <= 32'Hfffffffc;
7972: data <= 32'Hfffffffc;
7973: data <= 32'Hfffffffb;
7974: data <= 32'H00000002;
7975: data <= 32'Hffffffff;
7976: data <= 32'Hfffffffd;
7977: data <= 32'H00000002;
7978: data <= 32'H00000000;
7979: data <= 32'H00000001;
7980: data <= 32'H00000002;
7981: data <= 32'H00000000;
7982: data <= 32'H00000002;
7983: data <= 32'H00000007;
7984: data <= 32'H00000003;
7985: data <= 32'H00000003;
7986: data <= 32'H00000005;
7987: data <= 32'H00000002;
7988: data <= 32'H00000002;
7989: data <= 32'H00000005;
7990: data <= 32'H00000002;
7991: data <= 32'H00000001;
7992: data <= 32'H00000000;
7993: data <= 32'Hffffffff;
7994: data <= 32'Hfffffffe;
7995: data <= 32'H00000001;
7996: data <= 32'H00000001;
7997: data <= 32'Hffffffff;
7998: data <= 32'Hffffffff;
7999: data <= 32'Hfffffffe;
8000: data <= 32'Hfffffffe;
8001: data <= 32'Hffffffff;
8002: data <= 32'Hfffffffd;
8003: data <= 32'Hfffffffd;
8004: data <= 32'Hfffffffb;
8005: data <= 32'Hfffffffe;
8006: data <= 32'Hfffffffb;
8007: data <= 32'Hfffffffb;
8008: data <= 32'Hfffffffd;
8009: data <= 32'Hfffffffa;
8010: data <= 32'Hfffffffa;
8011: data <= 32'Hfffffffa;
8012: data <= 32'Hfffffffb;
8013: data <= 32'Hfffffff7;
8014: data <= 32'Hfffffffa;
8015: data <= 32'Hfffffff8;
8016: data <= 32'Hfffffff6;
8017: data <= 32'Hfffffff4;
8018: data <= 32'Hfffffff4;
8019: data <= 32'Hfffffff3;
8020: data <= 32'Hfffffff0;
8021: data <= 32'Hfffffff1;
8022: data <= 32'Hfffffff5;
8023: data <= 32'Hfffffff5;
8024: data <= 32'Hfffffffd;
8025: data <= 32'H00000003;
8026: data <= 32'H0000000b;
8027: data <= 32'H0000000c;
8028: data <= 32'H0000000d;
8029: data <= 32'H00000009;
8030: data <= 32'H00000009;
8031: data <= 32'H0000000a;
8032: data <= 32'H00000009;
8033: data <= 32'H00000006;
8034: data <= 32'H00000003;
8035: data <= 32'H00000004;
8036: data <= 32'H00000000;
8037: data <= 32'H00000000;
8038: data <= 32'H00000001;
8039: data <= 32'H00000001;
8040: data <= 32'Hfffffffd;
8041: data <= 32'Hfffffffe;
8042: data <= 32'Hfffffffa;
8043: data <= 32'Hfffffffc;
8044: data <= 32'Hfffffffb;
8045: data <= 32'Hfffffff9;
8046: data <= 32'Hfffffff7;
8047: data <= 32'Hfffffff7;
8048: data <= 32'Hfffffff7;
8049: data <= 32'Hfffffff9;
8050: data <= 32'Hfffffffb;
8051: data <= 32'Hfffffffd;
8052: data <= 32'Hfffffffe;
8053: data <= 32'Hfffffffd;
8054: data <= 32'H00000003;
8055: data <= 32'Hffffffff;
8056: data <= 32'H00000003;
8057: data <= 32'H00000008;
8058: data <= 32'H00000006;
8059: data <= 32'H00000008;
8060: data <= 32'H00000009;
8061: data <= 32'H00000007;
8062: data <= 32'H00000009;
8063: data <= 32'H0000000d;
8064: data <= 32'H0000000e;
8065: data <= 32'Hfffffffd;
8066: data <= 32'Hfffffff6;
8067: data <= 32'Hfffffff2;
8068: data <= 32'Hfffffff6;
8069: data <= 32'Hffffffef;
8070: data <= 32'Hffffffee;
8071: data <= 32'Hfffffff3;
8072: data <= 32'Hfffffff3;
8073: data <= 32'Hffffffef;
8074: data <= 32'Hfffffff5;
8075: data <= 32'Hfffffff7;
8076: data <= 32'Hfffffff8;
8077: data <= 32'Hfffffffa;
8078: data <= 32'Hfffffffe;
8079: data <= 32'Hfffffffd;
8080: data <= 32'Hffffffff;
8081: data <= 32'Hfffffffe;
8082: data <= 32'Hfffffffd;
8083: data <= 32'Hfffffffe;
8084: data <= 32'Hfffffffb;
8085: data <= 32'Hfffffffd;
8086: data <= 32'Hfffffffb;
8087: data <= 32'Hfffffffe;
8088: data <= 32'Hfffffffc;
8089: data <= 32'Hfffffffe;
8090: data <= 32'H00000000;
8091: data <= 32'H00000000;
8092: data <= 32'H00000001;
8093: data <= 32'H00000000;
8094: data <= 32'H00000000;
8095: data <= 32'H00000000;
8096: data <= 32'H00000000;
8097: data <= 32'H00000004;
8098: data <= 32'H00000000;
8099: data <= 32'H00000000;
8100: data <= 32'H00000000;
8101: data <= 32'H00000000;
8102: data <= 32'H00000002;
8103: data <= 32'H00000002;
8104: data <= 32'H00000004;
8105: data <= 32'H00000002;
8106: data <= 32'H00000006;
8107: data <= 32'H00000006;
8108: data <= 32'H00000004;
8109: data <= 32'H00000006;
8110: data <= 32'H00000004;
8111: data <= 32'H00000005;
8112: data <= 32'H00000004;
8113: data <= 32'H00000004;
8114: data <= 32'H00000005;
8115: data <= 32'H00000005;
8116: data <= 32'H00000004;
8117: data <= 32'H00000007;
8118: data <= 32'H00000005;
8119: data <= 32'H00000003;
8120: data <= 32'H00000006;
8121: data <= 32'H00000003;
8122: data <= 32'H00000006;
8123: data <= 32'H00000004;
8124: data <= 32'H00000006;
8125: data <= 32'H00000004;
8126: data <= 32'H00000002;
8127: data <= 32'H00000004;
8128: data <= 32'H00000001;
8129: data <= 32'H00000003;
8130: data <= 32'H00000004;
8131: data <= 32'H00000004;
8132: data <= 32'H00000002;
8133: data <= 32'H00000004;
8134: data <= 32'H00000003;
8135: data <= 32'H00000005;
8136: data <= 32'H00000003;
8137: data <= 32'H00000002;
8138: data <= 32'H00000001;
8139: data <= 32'H00000002;
8140: data <= 32'Hffffffff;
8141: data <= 32'H00000002;
8142: data <= 32'Hfffffffd;
8143: data <= 32'Hfffffffa;
8144: data <= 32'Hfffffffc;
8145: data <= 32'Hfffffff5;
8146: data <= 32'Hfffffff9;
8147: data <= 32'Hfffffff3;
8148: data <= 32'Hfffffff0;
8149: data <= 32'Hfffffff4;
8150: data <= 32'Hfffffff7;
8151: data <= 32'Hfffffff7;
8152: data <= 32'Hfffffffe;
8153: data <= 32'H00000007;
8154: data <= 32'H0000000d;
8155: data <= 32'H00000010;
8156: data <= 32'H00000011;
8157: data <= 32'H0000000d;
8158: data <= 32'H0000000e;
8159: data <= 32'H0000000b;
8160: data <= 32'H0000000a;
8161: data <= 32'H00000007;
8162: data <= 32'H00000008;
8163: data <= 32'H00000003;
8164: data <= 32'H00000003;
8165: data <= 32'H00000001;
8166: data <= 32'Hfffffffd;
8167: data <= 32'Hfffffffd;
8168: data <= 32'Hfffffffe;
8169: data <= 32'Hfffffff8;
8170: data <= 32'Hfffffff7;
8171: data <= 32'Hfffffffc;
8172: data <= 32'Hfffffff7;
8173: data <= 32'Hfffffff9;
8174: data <= 32'Hfffffff8;
8175: data <= 32'Hfffffff9;
8176: data <= 32'Hfffffffb;
8177: data <= 32'H00000000;
8178: data <= 32'H00000001;
8179: data <= 32'H00000000;
8180: data <= 32'H00000005;
8181: data <= 32'H00000004;
8182: data <= 32'H00000002;
8183: data <= 32'H00000005;
8184: data <= 32'H00000009;
8185: data <= 32'H00000008;
8186: data <= 32'H00000009;
8187: data <= 32'H0000000b;
8188: data <= 32'H0000000c;
8189: data <= 32'H0000000c;
8190: data <= 32'H0000000f;
8191: data <= 32'H00000011;
8192: data <= 32'H00000011;
default: data <= 32'd0;
endcase
endmodule
